��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d�
�����@Xk���Fq���$Z�u�չ���J 	��Ǐ�J;a��^��?�o{̛�����-6�]`D�F�XJr�ţ��ynJ�yj�2R���԰�#�P��>v�y.Ee �6�׷y{���iP��nz�]%�Cd��*�'�[������`����Ǟ�H� �a�C�����c�
|��iHO3J��U
la��h�N�'UӴL���e������A�Z6���.ƴ�3�قmb���P��m�x�:�Q��Z��r��O�Q>e�6!�G��`�V���
~��ȥ�!H��p��Wb�2���Tg�5�W�f�*L|�C���])��|�L=�$��ve�0�9���s4������d0e��pD��
m��yL��ߊ����F�q��I12��e�Hz���Ը1�vԍ�E��-iN{��J�#�|�O%*��\W�+G9�ثy�E(�$L��䜵�Q�YM��D�ϺCtS��h������SU0��i&XY�Z,�?
R����,�� �]����)^hּ�)]�?�@�I>�=l�[L:SF�+'�K�':��Jr�t��$ofu��g��pE�)�]�N�ep6�-�U�G��V�T�FrT�yn��͛�<>�L�_��b�D�a�3ܖ���
��: ���kOb���M ��� �w�'�_B/�n,&gz�Q�Q`�mJnU͵K���s�~�����C�KOe	s���^��m�Vb9m��=�g����}D�@6~J'�4�V�L�9��Z��s�)���)!䦟�O�>/�	#j�{6H6!�6���ˈ�X>��\�n� d�V�Zw� P�*�<[��5_�<4c��˝P�ح�v�߻�9��֤Δ��ul�j/g<�	��u�3��a�06�ߤG�D�0��֕��q�2��R6b�!�4��@Qi��rk����w|iJ�s��WdS�ދ���y����J���e�O�2 �Ո؇9�r�4����a�J]Z�f�p�Q�Ϧ��%���|'2i.�qv�����,o���C��R/5��[�$��3Mׅ���f
�z�7���T�_r
���wh�i=ǽ���Ao��S�`���~*���|.�4o�tX��ۘ��w蘑;>e��0�����Jĕ���� �j�P���zy�e�S��+��2��'�5�'|�h�~����%#;�gW�'��<�U����HN�����FVa����~���Ώ��m^J���_��O�����QT�֡�S�S�(��.f��9���`�,�{�1��XKتM�q�\�5.]��,Y�]���N�����RV&rn*`�Y�� ;���4�n�(�5���1~����p�E�-��=,���_K�?��c7�M��⁤�\}�����H��2S�2劖1��K� L��f��� �RAFu�o�����ͺj� {/��#r,��ǖ��֍�8Y�ۺ7Ld��,�3���Ať�]f����E�]���%������]�0vQ:s��k�<�4B8p��C���v�k;qgs�JT�3?=�%�iG��RL�Qϙ�h���|x��fQ�A�1z)�
�H\����F�d�;�.G��"a��N4Z~4���"����I�Nǩ�� q���~�@
�&K�ȣڶ�'^Û�\A�d�n�nt�o"�L�n��(U8�?�?��hw�TF-��DJVP���FT��$}�os��C6^�����}��(w�Ѝi~�J������},���5�sV���:�n��KO�%���2��/뙑�=x����S���Sk����	<�{�e�W��ҍ��o*�]l�1��쳆��H�-��ᒺ��i��=ڳ����J�˗��J��23�v�B����S����O�')��?[�C��Q^:�s(�}�z� ����r��^n:������V<��wo���^��"#��.,g�YD�ou��[YA�Q�d�fOJ���aA�/���:�:�~�!E�ӔK�L��^g��]%ԩ
������LML���GS���Â|&O�����H�NNsպZ����LjT� C��{��~T�.���� .%!�!�sW�jO�h\̣�;Ba͏��X%%�ʥ��p�%�'u����{19�!�O)��1�s���&<�G)}Ë ]��V����J�S�]-�u!=���s�s�����?�ŏ�"�э���4��iX>���R���9_v�t�b@����8��R!�k���0�TS�}$���Mc��AR*5�K���>����!�D��S���WZ��|"�*(�3{������u�iu:��A�{�dױ�/kLcW`Gt�	����t�2P����ڧ{N"����N���ʑ)�	�c\j"m2��ee��RN&�38��H���"4Su2�!j�����2�;���~`!����m�����+PD�)6g�0�}�Pf�F�E����L
����}%-�,qa��dw1�vt��Ǿ��{�x�%��ꀋ����v��A�-�Ax�o{zR����?�u�$_�߶�8*�_�8;tm?���'�0��W�Bs\����+n%خ�'���6!�:@����}Yxh*��{�Ve;*㌐$��̦�si^��B-R��TҞ��?b�������/����Ը� ��pQt�/W���;��7 Ժ�3m�^��9-�>�>����}���.7���)��m�V!�v�(#W�0'�y���"[��9�����HW�"a�cB�+뽀����b��h�ޓL�DV��9��A�|i��"A_���u��3�k,F�^8���t���g���`G�4�,���J�!JKR��1b�[T���I�D=F�L��q\����4Ͳ<�d�jX
p'�c���X�Ws	G�c��Z�A����X���<Oy�G)�5PP�r��㑑�uC�G�^�������0u?��!= �h���xV��ˤ�yn"��(O?4_�d�|нsͻc�+���T.lP�u���H�ȒtP!\���B��;����^���-�mߑ)�ha��#�X�;������i*T��C��+�'����W���� ��o�i3���A�Pn�K�4��(_-&��"s�gp���S�^Vر�\�� \�ѮB��y�_�>J��[ ��{��[n���t�gu�����:b��0����oQ��ٛ1�l0�|�kY�%rqg�@4hwL�=m<���u��lz��\��I\{�~q\2]cg>]�<c]�p�o�a=��-�t�k��3>�zL�=U:��鯇	@%��ubN�xWB�K�X���T��	Uu�?��O�l��$Ɣ�朩X��lI �W�=i��X݀㰲纪�� lN�)%��})��6��=��i˽}��(��ҳy��3;�oH��nފ���5��	�la��Z\�q?TjS~S.2T��)�Qs��bΤ
���~��j��H��&�ڻw/w#V��,jf�����w�(Q_kuQcFC���2/m�l@�,��_��6�0���;h4�j����j\]r+���q�t;��OUH)���6�vX�qVp���24�ײz�.'���s�U�\�1���3�Qan����ȣo������B�2��S300t�k�/W#sM#�e��$�B2B'+��K�ӣm��sZ�@Z)�]�FJ�87�zc��k������8�I]rTF4 ���ǓcZ���C���B���B[h�#�*c�D���Q�P[~tڰ���(g�{,}]�^I4UBR.%�bV/m�B��.�=�bDOI��#T�}�9�@\gT�]i�.m�8=2'
�/�BP���փV�.����MB�Da�EÂ���q�{B�/د���#-�R��4x)$���v���������S��Nב!�F��_vS��Pj�Ldpf�qW#�&�BQgD\#��.����՜�M��-l�F v�-A��@/F6�j��( �5��p����էx��3��i#�8
���.b�Al8,[Gב B̟pB�����h;Yxe�(�?4���f�����8�CH9�W����i��<��Z���7`&JB�U���z�A�������H�1�6�)��ֳ�z-�oE��;��XJ�ʙ>gM�C�T�"0�j�T��zmB��
�<�����������!�D�(�ƚm1Hn��A:E�s�� I���j��`��R�A��ARUV)��^��뀑�e�_N$�y�8̮�Lj�0e���:�F�.�H�j�T���0�ؑ�s��O��d��Y�.�{�6+�N�&�^��.i���Tjɹ�+�5�z7��y���0�sȖ��'#�x�Hd�<�-�%���8~{�\������p�x	a������!�Om�=��~a���B�3H�0Y��琭!��q:}�4&��b���%����g�w�3��kk�(4p�l�I�1]Qw(�Ar�퓘�s��[�<�~������ɭ
�"�y�Ї<�G���#<8>�$�#��#m7"��C��{�a�b�b�I�?�}����(I�E�Z��ӳ���΂%@��ԙ7��O%��-h����#�5�eQ���,2,�[ѩ����|���'&�7�?�"P!m����ܒ������E`M�tfc>�⼙�;�ۈ<��ҏ�;���}���3��b#1�!�P�8�kh�I*x��rU�ȍ�y������V��DE#O�?|�c�@��nt��lJ�pl��������'=8�{�/�By8	�$ZǓ�6,�Lا]�H#B
o6�2bl'η�u�C\+��i�h�Hd��V)�BάH���;p?��Ҩ�r��a��؄��}��{�� ��0v�
h?����a��}(t��Äuov�Y��77�뼚j<�1�d�T���t��(�K'Ph#]���,�}�v[yqG5rX�
��hj�V�Ki�҃�%�30bdP(�b���ׁ����	9��{"��h���#JZ�~�����	��T���>�K���>���'���UNY^����)�Q����.�p�Һ�8s�P��}C˅��Yb%��}�$]]�8�\<y���8�C�Wg�j�:d�	���̻~7R8�^�PT��-A�}c��KT�".��5��a���r���E�k���7b�I��X�GP���"ɩH
�f�d8^m��%���b���H"Q���d0Ɩ�� ��ʵ&���ȁ��b:�?dD���v2J��V�Z@��5��n\׭�>�x@��	��=u�3��z�����et�iE�j��b�~�S�4�G<��6�<x0�n5��&0żZ����cpS�"i�>��x:�k[�ݔ<�}u]�/���[�;�Ә0}�|(0�N�S�OsxS�����C��U���[�:u�GNл&,-���6;.�z;	N�4f�[%����rg�҅(�ý��B%���l���z���A�[�������*���G�a��]ZEIZ6��$��/�U��g�
 �����^��.rq�
9V2Y�=���l�{��3�fR��/�Z]H�y,�_��HR{c:�-��3���9#Ķ�&��&�~�4AO�A�����Y��D̳:D�z	��?S�@�!2��ol�x�Y.�w��`=�+���|yy�k�׳�g�奊�aa�X=P���=�&5xؚ�rf�X�>�����Z��F<�Gr�I}9`t��5K�;{<����C��
���p�&�*-k:=�s��).�;u�A��h�#jsw7���f7���+0z����'�@4�cPj]ϫ}G)�{"���p�Oߕϊ�DX�Y�Ck���]�o����!#s�%����;._ Љ�U�.@�Ę�<�����9�l*������|q?�T��S����;���TWy�_!#��q����H�&��[�
�*�sWK.�N� ���"a�����%%����f{k�6���2�H����Do�Ee���*�y2:�Q�9������^E��z�B�"��9	��.u&��O]Ü����C�	�W�9D
��'�Ý-��#wG�S��~q��q%0�p}�[��Я�����c\�6�oG��U��W��h��S=m+��_M>��F~�2=�q��}�l���.ʯ��"V[L���Z7z2][|'p�
	@�>�<�E���aN��ھ��r-�����Z����Xr# 4{�щE��J)_Aa���eJًe[?�]$Dv������D쌫!�C-V�blЕ��K�[�fǉn��̖(�(@�:'5��d:/���ߕ�ĸ�����>qQw�FB�!���ޗ�q��,�[�9z�.b�2�!�esi0���jB�pL(� Ĳq�K�+�t��o-�	%�璬�Z�IA�s^�+4�X���
���S��9������ۄ����g�6�"�i������5CbI�ˋ�	���ÄȆ�r��:F��)q�y�ң9����~�5JQ�nP��L�ash�=3��m[P�kt׊�Fv�D� e����K�6��4��P�|�&r朖��X�'@���B@t��V0M��*��ܬ�����wr���u��=Hp�E-���<��P6���T�Y�_C<v��!��c���x8s�SՊ�
w˭�%l�~,$�.�ڜ�::=k�8Q0��N��w[�����k��#�N��u+`̛Z�����v�6�%Ȩ�~�gV���C��W��		��} ��1f�o"4LJ���1�-F�e4�y�f�D�-`Ce�3@�ݽ����Ā��ar.�<�LB���Y_⇀ʸ���P����-�W�l���&�8u���m�%���Xunp��������&������\�终�����MOԻXۭv����9��uH$��Cx�����R�OKk� #RIX .����p�W���L�j9��ؼؿM�Dۿ��t�\ڔ�lO�W�.�t��'0%�a�'/^��>v�CLgFx��,Z�^�M�2'(�rP'�|?���ޮQ�0:��83�t|�b��O.�JF�'�t�&ݮ���|6�a�J�4hT�*�P6��Ė�jE�-�XƹLo��06Q?��f�O��a���&�^�r�����d��f.��K�{f���1w`��ٌ�y�ZUa��`���v\M�N��|�@�̫CDꔊ$'�1҂�[�U����g3�ĸ�K�T�f ����R�0�w�e��!9F��������\D������rK+���[�������}򿸰^�p\��_��B����(�H�����e7�Q����7Ɇ��I���y #��+(�������������t[+��R��Z�������zE�~�v��Q��<(LЂ�|���R�>䃞�8#���`��/���)�@�i�M�GP&۱��E�Q#yҩ��f�{�-��Cۘ�ٛ�K#�=y2y�LGԐU�
�N�q��:[�]wg������*Y/�����x$�L��	�5#��?w���~u1����Fj� H�N���-� ��v��?)�"��3�5P����#}yhG��%rX^.{�C"�2]h��s��W�/&�U.��_��|=p%ݞ�p�fv�th���<��ށ�N��a�<:V1>�,�}����9 ��R���$�n�7CSR����*[uv͌m�H�w:+4D�n���*��ؖ슉L�1ů�������r�QV%���#T&�*���6P��F��3�{(�lWޠL�t]Ù�����rp��8�=��<����yh��)�)qa������j��Gd`�&�`�&o���� g�%x��Q�}�]� 
Dt�Oo�@�_�bi?�MW�����f�$�q���%�0թ���K�N$����Jmdd.�ݱ�=�Ŏ&��19s��Nv霮3��Lo��'�� �&sh�e`>��J1�����*�z˙�TzT)�M�Dj�]��K����cig;2�`ôC�y��X�����Y#��'S9��I(���X�Wtt>�v�J�F�A%��|*�u���M�u�p�O�tV�v�D�6�̇
{��"���]��V���킂,0)���0ڡ�HLWOe3��$ޫtPRug�Gn�����-�����i��u@ܡ2�aB�ªF�\�$����w��=��{�sZ�z3�13Ϛ!5;�<`6D��.�F(3�J�b��
���SE,�iĆxK��`��M���r{�IG!U&��a��X�u�<ustj�>�2>Y�e���g�p��-:;.��3��2�d�7Πݑo��y��y�%i�d���ߒ�J������-xm3Ͱr}\<8�a_�k�5:�3������om&���u�xȇ���d�?`���lVj������2�i/�Q��)��?_�[���Kt����Ӭ�f�����W���x��,:�������F
RI�S}"v]1N�wF�z ՊB�zs���MHc(�k[�Eh�G�L���-��}��A?�����Jj�4��c�O�WrW�Ӝ�����d�"}=B_,l�l���^��31�UxϞ�$V�)x8+�DӅ�F���_��3zK<^���i�k����V�B;��������w��|�)�:��0Y 6ʈ�l<]E\��s��\B`�!�MB�S}5@Y��%�O?�T�Sa�|�*�DzCs�R�/Tҽ���8� R�5�AL4@�, ?g�iQ!����ǽ/�-`�|^{c�^�p�6�eR��<��a�w��xMgJ��n��T�xh�
���n�B�\D08B�Գ.@��Ӽo_��"Veb����y[��~8wA�Ḃ�F�Z�SM�y`��v�����P��7G-G	���964{��@%�[��h�� ;��[�L!�Nh��j���Éj[$�6d�Bǎ5�qAc���t~��y�7����*u�X׶��=G;ʎ���z�����3�����a�����V:���f�^|�E�Hb�V}?d,��0{w�`��d���	�5[��qp];X�� u��swb��.)� �n߱1|�\�`�!���ц*+���z�������d�	�ȡ"q�ה�<�  x�~����y5	B`�L2��r���<bA�JJ�c4;�xI�'��~����^���e��|��ͺ��tJ *������z�"�b��X��?!���͢� KE��%p�^���y����k��L��$h����b]-E
�w�an���Bv%c�]�*����5�CW����;/w#�hIg����=v��i�Α.\��k���l"���4��t��|?�;;��nlM�����Q�6��,8T��\?��
�������-�� r�z��`��./ ,�h�W׋� @��A�<���ΔI&�&��x�?T?7~ļ�R97�( S�� �v<���Ϭ̔)��:�.�PrX!�u�'	�y�LG~��^s�6*=$V�W�_Ѵi��t��k;TvP��I�%�زLMX�\E�U��y}CB%�s���������>t(ۢ@)���BgR�����:􉶫�֏�	4��ghLxx17�Fї���_t�[�Q�;aL<`��fk`CJ�P88._��ؠ�3d��b�W����R��'���b�q�~��h��T��=::��mp�.�q���0�������}Oe���?MN4ݸŌ��7p_�<%$Q���Zz�E�|J��ħk�#���klO
k�[��(�]#��ڗqN{*��{�{Q�1�L��6y��c?̫� �KG|�<�Ҝ����������W�a�H�>�����3s�6Ÿ*��a���_x��R��+����z&k����ڎ$�D1�ғ�w�`���B��5r/�?��_XiKy�%E��g�V���k��X�מ}c��y�0��)�:�Tj�v����Jç̻,��;з�	}���O����9���no�.��8�o�[�O��R\Kj�0�*�}�����N}��=�o|*P3��|�c�lS����L12�e���Mm�+>T�D��\�5n]j4��i<<{=�]�߱�����9Y�}0��UN�Ѱ�tiv���#��;-S�׻�7�X>� t̎�K%
��P����`.U"O�٭��j��ݮ��oI�Ope��sB9u\�o�k4i��La�t���:G�����Dqk��5�� ���f����Z�JnM]�$R��V�({<ݦGa���rqȥpq���Nt}�_�*$<�SF �Z�%�יd�-�������x����,�@A�3�<i�GGhR�تC�l\LԌ�ԕ<i��X�Y0�CA�J���x�P��YJ��oH2����):�� `aA�$=%[Ԋ�AT���dl��}W��n,q�����C~�_�_L������x�H�J�Y�_��#��4�5�:p�;�ɧ�&��*���a�1S��'����<!x�F1�,��@�{T�`��{´����,,�\�رO>|�m(�%M�m)����7)�sl�_Q���#VL���
H�@m7�$Sm$����>�$��RE�n¬2
�2[��T�%
U��g�eL�X����n��O'��Y	��P}&�T7I�6���~�sSWhq�����U �⛈;P� NS�H̷��?C��=QPu��u�P����-P�{(�]�Lw�<�(E��x��g\͆�)\9�:FI���}�ҷ��r�*s�����5Q8i�ʀ��NY#K�E������0�\�kz�Y���#D���)l2Fa��nc޷��?-H�J�@�,���se�_��
>������H�E��`[F#��^�L������i��\<�� �̞�E��L:���D�vRv�^l�@nА��I1����y^61����v���
����_� P�B��]�LjҍYp��<8(�>�D=���"���#��`r����eMv��&�w�0dUQ�ST�`���2����d=�bK��ųTW��{�����u$���LmbG�ħ�i�IILH�8�B�V�N�m���mQ�?�Z�؂O���+M3\m@4���nr� Y��#_`m#�j��ή�!�����Aak��]/؋�N�����E��6�=�n�D5 0W������c�0��[s�%;%�g�����z][�S��g��f�§Ɔʯ/g�s�6j'��K�=R���
Bv���\�y�h�s�О�U��F]KB�`x�NALzAv|W��@��dGe����X���̈́Y��!�>/�f�mr��5�?��>��9�f�5Ġ�|���xk�$����(>熝j1�*묟i#���
׉oߗZ�i���Q�wf=l�nw���������|L:�'��":נ�{��xaG����X�_�	������3���L�lD���H���f[݄0J�]#PPqKOc�����P��Q^Խ[��]��%o1i��ڤS�Ev;!Q?( ؀MVN�6�-{���������:�
:L��j�Ǟ�7`���3�H[[���WB^�d���
8�H��f~jkXig��{Ɛ�e+pnȃ����ꑔ��SdϠ{���K�z[�=S��d�Ͷ�(��6��MN��%�����jw��O@��,f�����@��V�%	7�����D{�g<,�N�u]ORcey7��2׭� �a;mu����c>�65���蕓��d��oP��@�U"���Hj�J�9��c4g�]K>���$v.���C��Y�fF%&i/�6�U����� dX.�g����Czk�>�&��FZ��xqd3���,�uN��8�g�dW���k�>ʂ����S���z�sk�Ɔ��Y�z*ǚ��_�Z7;		W��|�mnS���H��)�9F��$p�i������3�q���4�?�|(JK
ЬHը����@VY�D����"Y_?7���XѕV3�K�!��y�qNW�F���o
ZFPh�I�� �q2�2�V\��q��s6�z���R�'Xj�������iN.A��6Ye��_�㕩�=��[�%,A��P/v�eT�?��ɓ��O��}h{K��� �s���V]cʧ�XP���r�� �� \Ts�ļJ)�����릏{�í%������#Z�09iIMH�f��q�� �QZ�d�&V"�1���L�!����]���su�d��Ǧ���5��f�6~^��~:�����6F�5�n|�<)0Ce�L�&��0���Q�+󭍏;S�>�W�_H�'�ٰ�5��N�3#�w�!��X{��|F�J�kָ��Nŉ���⑥�㝨�O���Б��5�ϯ-�~��Xunɺ�2�2+E9I�j��Ҭ�g�P�Hz9��:�ER@�]aL�M���JD��åZ+�Z�+�3_��R���޲>�d�N=9!�'7T�M�Ļ�����c활Q��8�9�6;۞p���#�J�r)��'�vR����y:5%r���J�Y?z"��H�#�G��p����/��tT#K1]ˌ9��p�Lw��ȇS�@n��e'�-y�CF�y͓�'���셒l�6���f��`|�ҬEEf嬯O����i� gQ .k>���ˈ�^�Ϻ�!�¿d��p��gf�
�q9��w0x��"��k����l��`���˕���g�=�vY�A�)�);V�dQ
A/̥�����2�.��3(��]�>ڱ�~�_/�O	um�Cvͧ0�d�$M�]1oӲsN�u�I,Nd缌�xQF����>K��>&�$W�%��9)��\d�%|?I�N4��dI���R�:^��hb���,�/��X3i�m}����ہ��7�E��s{l�J��J͊/p��)���`�W����rg��0V.rp*XB�wؐ��44?��8��
�K���ֹM'p"�Y���V*׉e�9���ʏ�,bY����<{
�&����u#�J��iS>9Y|������N��A`��� Wiq	��˔wr�.*���~�r���"Kl�
��o_����wY�	�oŗ�WP9A��v��,	��,Mɤ���HjAD=#��q5i��t?�^���q�z��;�1m�`3�? q��fhg=j�ݽ!Ie7��P���<7�*�b���q����9�̹A�j�1�����8LH[�>P>:�~�o�yFݹ�y$�N��Um������'��Z��Qa>>�5/	�g�`���K��[Q�!lW��/���hW.Ws�]���Yd�^�@�ɰ���Z��a�:T��=!F�B.�W��84x��$=?��bZF=Q�o��&kXU�,��q"��ek�RqDPxm��n��25�bW�QmY�3r��y(z �Mf5e�Ή�r�V�xU�R��ۥ�1��ƙFc���U�A��&+�V�W�ˏ>u�בȔ�rx'�:�[��K��RA%V��K���P�we���l�f��q���9�9��[p�͙>�gm�0cP���^��YI�2؍$J���x�B�T̖���i��%*�,�P��<��0\�
�Ӣ����8@JI��7��^�i�M�_1�J��9n&�T�^-ZL�=�If;�L���s������D��{���Z����Տ���@�����`���h"����ߚ>w �yB3x{z{Dr�rY�3��ƣr�&�b��m�	���f�p��I�:��M?i��~q[ۣ�h���#�;w[�W�Qͦ�'�X����x̽��e��e!��
�f�_��qkG[�'�BM˾���鎷W�9�A�1�,�2J�\��W�i��#=�>Z���N��x�a��-�H֩��P�ȭ4�}5��(�A����ֶ�Y��譣�8^"���^��&ס���;��4�x��H6�b�g��l��q�7�m��WBMD���8�������g)�C�Z�'4��0�0t牌v��F�����;[H����B~U����&[����c9,-$F`��R���bj)BE�l_>��5��^���?�sR�8M�;��� ��ر	�i6��G甤�#���/�`���@�+�L�Ѝ�[C���Gd���ɺЕ�iF��7$ٟV0�@��T.w)S53j��@"��4�PRp�Z	�Ƌ���#�$�W�K��⚌���j�c1[���h�1�|Yc�Ff:�1���}��h{}�}2���gf��o�a��!WJ����׬Z^���9�s?,8��d������L��2h����"��F�Ʃ����/�s�vw2�U	�#��q���¤�
Ғ��N�grr^n�X��Bg��*j�A!!�h!���n�% �~�� ���O�I�h
L�!���i�hT��������FO}3� ��@����� mɺm���H����ң �(#R{㷬�ywH�1Og��l;Ap_aS��!��R줣�E4Hxb�ث��bv��������/�\�M${2��Y�~���b�5(��HwB�Òd��H�k���	}-:���D�)��o�I9��"����1V���.\�j[-\��\3��Jg�X��1�F��~UZ?s��ɤ�  �ae�R�`�z�] �Z�3��Q��%0�Π�K9�J���# )U*�C�#F� %�\��!ێi9�&�$��<����*z�L`�<G�k��'-\׿mr��Ѡ΢ձ���/I��ۼq1���ޘσm	��)�X Z;�?���yϛ@睍�)k��[��w/���5�����;�?5��kV#��ԏ���Y
�>յ	�^�-��]��W݊9ƀ �ᦝ͂�6K�2��${[q$xk��g�����)�*,d�s���J=|�Њy	�E6�):�E�R*_R��d�e�������Q�pX����g�F�	�2YR�Ǹ������ke0��B@�Y�����hs�x�"�����4��� {��^����.�T^<��h�4I�|����T���P^!�pբs�Ra�O1W�?����n�;��n�	�����$�rC���&�F����\��t�^�N�
�O ��a ��5H�r29�Ժh�����J;�ŝ����]Vє(t3:ZmzY:l���R�,��mߕ+�U�{9O��Y��B��	DaW���X��h��}�"�Q�#g������Y�d��2rF�
���-$��?����Nl�!�p�?8�E;����qJV#%�����a�N^��������f��\�kI��t=�Y��qᾘ,���g��!�8�K��:+�/���t(�t}:�T7d���ƻ�/K�6Lp��({����f��Y��U���t�)�}�����х�k�����4���������R�:�kq���K���Fe^M���ܔ�ey�a�n���WPp�\����C},�9}�ή��.��ָ��� Bq�0!�{D`�Y����*$'U��5��K����+ִkU۫���1C�]e���Ś���t�� ���/PAv @��t�U�GY0�$"�������@�kP���akfG���FXu��<]�6p[A�x��Ɗ�b��bˇ�B�@A�D�BQo���bfA=ZL���'Y@��p�>�P`63I*W�W(�{�\��5�|k[�~!㢚E���p7��1&a������PlW�?^�0�Zj�G�eg�W������A�����ܫ����-¢z���e����|���<��r��Xj�yq4��K��s�_L��_�6U���Q���V>�f��~�6Xk�,�T�.R�>`�J�Eг�hFpyI� �Şh<Y���"��� �r���E���ʊg�O�s�[�F�>g��-�S~;�- �����f�4��Γe yp��;^ ��Ĩ� ��c�� -��pP�»^���^b5���Q3tlpw�N}7K�j(d�^0�ܩ��yr��tU����4���h��0/wb���^�� ��:�I�h�}�O��Z�>%���_P�A=��^kȮ�0h�&������%Y��]��Z�]��i��R��Y���ᦼ������B�"�1Q�����CW֌��h�Tu-��l��L�4e�c��p�AyˎX�����qI%fƍ<坶+��[��Ǽ퐾e���'[]�����O&�k�H��#	Ĭl��1���H������B��`Tj�&��U���ox���i|~�F��t!K�������U�WY���/�g#�@�Bi� 	I�vs��9�����u���3��>��� �.��|Y��mh��t����u_��٨�%��y��>M&��RY�I��+�m��+2�����{��Wkls���u�,��nЖj0���k���\�����g��=��[~�z��j���x��4�m�h�q�̛�;�=H�k��<s�o�$�yW��)$81Ϝ��Y��u�*��^�^
-�{�4��T8ߎ-�������}��ی(#Mi�K�P'h�J���{���c�!�񿈌�=�X�����뮽�Ka���Kh��f��RɤCl����Y����|<�����|��%iMSy<p��';}e'�ԁ;ƕ����a]���s�/^&e�y��,��U�y���m��q�H�ༀ-��כr*jL�3o����	4^�!v�"��+�WG�����XtG%ͻ!��N�S�p�^�nd�Ô7C��l�6��bI����ihF�%�}4f�r]�MZ�6���j��;�G��
{ ��N�-e��:b
wl�B��D_�w_ؓ�ߠ%N`���d{"�U��h���w�[�8l�4\j�}~�UN.ڦG6��,]����++hj9���k�z���F�e-7���s�1�ڲ�)K�_9\a��ᕤ��)��:<��s�\~��5���2G,�v�.e\�сj O�����	�X�S��`6���$$�x��1�v�8�����&;��Mb.'f`<�����L���g��+���ω�W�0����/��ˇ���UP��>^��q��
�ubc��������fxz���!Vi���N?}��&�!�;�����u�@:��P"���`��6��9��+��V�Z��l���2'�|��X�wL݄,0`�O,S�u[f�qGnE���4�
�
P�IjY�2���D>�L�ϯ���>��P�A�<��
����h[��V ��K�T���[jif��N �0�Nx�1�}�sz�|އ
�mg-�(l�#��,�F�*ρ�Ψ����˘>w���q�F�g�r��������d����BAAEx�������h�V��J*��]���:�%RC�2l��D�5��(n��kl�[5�idHm���Ή��4�J[Ȗ���)xGz���L����ni@����ɵ���4/���Hׁ�"�(I����mO�{E���Uz�2\6J���Xe�6�	��]����>尰����C�c�R�}J�@$@)���y��/���jx�'JM����af�LU}��Foc�8�I�a��3E7�O�1����gv8$����ђP?_�9�_H)Q�N*��/��j��_�a�F"`�a s����g�	=���:B��~Rmfh
&4
�5 =��7�έ���C��f1����rwx�ʑ��1 �K7��h���@��9�O{�2����y�V,t�FK$,\4�{!�4��	�μĀ��3݈[���_�/�yҚ;�;ܢJ��m����_����<$�se9/�W��L��'��,_�׳�^-kir�I�L��Q�݄�3|��������0Fٜ"�Ds���hθ0���$��ȥ%u%g#�^j�vʧ�4N�.E�7��U6���o�jd��v�=��1�;��%s�)*�hV���|Ui��"�~�>�����B���!�e�k,�(�6a7���������|2l�iಸ_�A���YBeWpE"z�Ū�G���z��	�9Y�r�hB9�t)�އO��V m�t�Ȳ8�c%=��:L.��[�к�6'���|���]��IB(5DOY\���.ײ��d/�0y�d���N��C��5T�Ӎ�g���s�< R㫔�?=�v��E��+E�m��[�?F]#��k'l�O��)F-
�����vh��V��q�Ï���3���W��.KE[$�*�����]�!��&�M����{ǝ�4��J��y�}f��6�E�/��ň"\#.f4�7��r����Ƞ��b���ױ{w���V�Z{�Ēb)n0&u�$JE=$b
3����І�f���d��(���,QгJop�k��2ƙ�K:Z��z2��2����<��s��Cb����޸��_�^��&��%�b�-Ac#������y:'���;�}�Uڠ	��DD� �<2�y�lSe����9��(�5����U����xJMP���^Iz�T��U�;	#�Ʋ�xN���6�\�x�w��~8�\�6#�L�x���,�
�>�S�y���x+���ݟ` c�r�Y7w;	5��a����r�"�߷��~�[����\'��M
t�G���za�z�q����
�"*T	,YNz�(� DM5��?+W3zM�2�����T�89s��	�:�П֮)�޲����{qH=ɩ��,��P���n�AޮE��)�|�
0��c�?1	��j}ǉ?�̐ъ�gB�hN"u"�~��yD�a��u1�]�V�_��g�Vs�ZF��H�'���r =i+�����2
Dq��|�˭�2�F��u��aIr�j���YQ*��K�A�S-�3�w�Z��m�����r$�}�T�op��T *Q�+`�����ߥT,"E��fi��%P�O]Y���� \~W*���1&7�A�_![��.�o�8[�o�s�'ײ�qJ,��7*���]��s8��2�s��S2�CI�I��jw���ub�3D����+���,N
�iKցjr�NG��(.�p��3����l^O5��/�_����P;i�V3z���n��Y.���E�����tX�nA�0��O�^��$����x�˛2�ݷٶ��A��H�=�S��(6�#����ASD�}��+^��>�坁ʩ�^������l��H<�f������ԭ�e��B��k.�SͰ?3��!�:�K���4�Ɋ3C[0�q_-e \��e|~G�y� �e9��=8�3�!:���K�r�;C�+Z����g����Д�
u6݌��R���$�gU���>��S�]9+A%	/�:W�X��
d"&�l@`i�'jŮ�]6��.�[�f�K��o�@S�gfϲ�;.i�?X@K��r9	#
.�EJ��`XQr:��=�Q" %�7��5Uʳ���XD��tȚ�#b[�0�-O����r���l(���+�y��\���qbP-@M�������b4},�?kVe�2>��R��(�*�.5��T�Ç�y��f�2�F�S�W����J���=���� �w"q���� �֤7�W�����Oz�,D��^B��v�A��(Q���Z�DDEO8i~kH��MBd�(��/����'3�$��v��kq�[�EQ��ܽ��1�����%.�/K��� ��jD�\��]��쐄��^�>�6�U6z�d��ޓh�aX�T*�yW6�·ɖ���iX�T��������Oa��A"?QRq)B0-�L�V&U&{�	���VǠD>S0f�1ɴ-�Ϻ�
�~��/�/.���<�.�b����|�`��7X�E%�!�-䟃��O,;`�}$��m8����D����*��s�G�T�d��bM���B8�&�Pgj�����,i����������*M���MK�{Ǭ���b���-�?�j�0����GM��ǣ�W�3$l��%Awܾ�2�,n2j��b%/�Z�h�����Xbj�A74c쳇�%"ا�߰]ͽ.1���@|�[��P���?�$oa�@	��s��}-�-�� s����^�)��[V9�D���d��&�@^�Ip�Q�ԫ�*�~,S1���bc�XrR�����w��fse�!�~��� ��{)�*��ga;x�F�D�2��LT���r�]t���׹b�O8�w=s�1K'���$���ߣ���3���{����M'$P'�;%������� {eu5�:옛ĉ�"���F^���1|��`�۽*N�p�tO��X�󁓓�au���뷲c@3��i��(�Ɩ��=���Dɜ�'U{��#0�[Î���G�n�cɍ!	G��H(p��X	Y�~L?W��v��82T�M��n4�� ����S"��-)20#?=j��*�L�����h��V�*�nN�Հ�εd�ʬq�1��؈Q�$�;n�Mc�{m�x�R��x�Q���Bڜ�� 	b�(�m�>ƿ�S���v�U�-W�]w����]y�D��p�ѷ5���G:H<Na�ijH��/6����4��5���C�8�Ѩm���b(;����lu��@g}�a�/"���ۺ�>+m(r�S��� ���)j��X|��(��|ֶ٩�/�ӏ�]ӱ���$��ь&�-��O���#!`Sl�WY�(B.9����:��y�N����h�.�!�׻�}����yNɎ�8hX��l����_�����	�&ok���\�N�'E�yAd[��ɕE
�����އ�cj��0o�W�] �e\�3O�-���1�OT��I6�%��jHh.�Jg??�4@�gq �6�%R}ђp�F���ԑ]���2I�����@5'��g�W!Q�T÷�~�T���(�NJ���z����#ǣ��� E�̺d ��~�e2���`�$m
Y�N�_vܱfh�?®׵wآ&M�3���'GB�#3�]3�02��?���2A� ��b����x�'s��i��6�=���(��@��T���2w=$�l��c��Ǎ<ξG�a����N.(dʒMt��26��C�`�F�D~i����z�%Vg��������.�gL)a��-Z�S��޿�Gh�$�';^�|v�LR�]�)� ʠܩ1��W*���4 �iٴ��\�� =��>�g4{w�Y�H.��������z�Ì���/�ݣf �RS��,g>�����-z��]�4kҹ�fJa:\�1H� �2��9q�(-yS��י`붊l$a�[�|���e�UbQp�4��^6�y��:i���2���u](��-}����pΓ�pɤ�H���M'!1�$�Z�/X���D�7���k�;t�\Yd�^Q*&g��C�.\f=��R[�6)9�Բg1�x���˄&]�����Q���D ֕����Z̜̥�U�q�R(��[��,G�(����i]��\	�&"�4��)����f�/�a�Z#F24���e����]!�U�	91>�}�1Bc�޵p��s#C��F�Q�(��R$��L���9bc4���+U%���SPH�~�u����% �"2�+ �w�|d����s��`۬��1A�㾾���]����m����"���@C>u�c���[1b�)����5������餤�u�ba� ��e�����0�����l������7�#��eD��D�GX�﫶D=Ƕ����/Vv�h������j�������d�bl�0yzڋL@2�@ӑE��u��;f����N�!Jc�(,,�oj�$����Z�4(2�-��wӼ��9X,x+��nqӋw��l���+*�I�+��O*.}��d��ݩ�;��W�=R��I/��1�N�K`�e,(�[�t��qqVL��k�ȟ^� +�j��e��T�Z֏�����l�hH$��Ԕ��_���<��
�u���77��m��Ȫ䦳:����|Q������B��¤�_5���Kr4#�!tK��u�?�G\�Ҵ:"�f�����{(��q1`��?R���p�������h6��i�ܝ�	�c}h���ѥ�|!�����t���w�Kp��n�[�ڐb�ی�z�!��@���d�.[�딂���]���gݸ~�E�����c&:�@�φ1�9p�%����
�,*t/ZKsAc�;�"6���|�4��H���o	�[���"����<�d���������Wl>^���׋��܀��I��v�v�=�l:�l裧�	ք���������s=���s`�5�@1#��E+h�e/�'�� $B��Ք'�!Y|7�|�3��D��o�����?4��"�k"B^�:<��h�������7ʇ*3V�!����B�C����*�*#�;-Xp�(�3A|M}�����C�l��❈}�w��;�>)��4<����k����kL!��e��k��8�֭��֫����Ft׏U� �ٲ�GD���-�+@��C�0�/�XlX~#�
e=�����ZJѸ,������^��$G*�hHe�NlWhg
�����\c�����!�Y�l�2��,�gf�s�} ��U3����l��{�T��V� ]R���AD��-t���v�N��[�ݥ8pk��㫮0Jz��C�5��0�%�l�6@S{{��;�٣@S�,��xX�\7�#k�f���ǜ����v���R�� ���;U���6�y+탙{�5�2���,��Oђ=��������p�uA�A�i��-��t�.+��4� yzө7�w�G�����B؟�CW-�u�m�f*��w�Qְ��[��d�&�E�JxH��U�|h�Wg�9d�$K��� ��r���G�%�?��K�F��YʕcF�7��"c�ZA	ߗ�L�/F=ukYU�XX�C->@�SuH�g�آY5�=�ibB�BGdyB���%!dD9�wc�8�X�/ 0ET˾<?�?	>���r]�+I�xN�S�&�SX��;�E(@h�����v��y����-�E�3���FT���4�>m�6�kI��9�/p>K�"������ M�)4{�m�K{v���\E���B:$�����U���pV`�tn�a��q0��$/���%��Fu� 2��Bv�N��- �NCm��B�!�}T�j(�#�L� �9���!���C�jO��Y�������_��'��p;UA�<+X �w��˸�g6�-z�UASy;��@�zL���'k�;��U$oh�d��@��T� ���D�����]�"}��� �7@ȁ�-^��l+�XF8�b�(:��ًɒ/�u�y��ck�sy��=y�,!��s�A�P�V��Ro�L�b��Kz�ț��mT����]�����VP��<>31	�N�pp������]pZ��X�
��ܗ|W�-֧<[ٶ��'��NT��`��5+�4�� D����Iv ��W`�Ƞ�Ѫ����@ܖ��3��Kd�b����F�X�vT�%r��:W���RK}b���Uc�c �� �:�m���'���_6��P�_e��ӭR��}g�9&ܵ�Вm��1DD���5[F�"p�pW�)�����!T����� �A��.u�=�y�n8߉W�����TX�>Wv�ɷ�8�kW<��s8����QW�<�å|�J�Q�[��-��g}�q�'�3)V�2��Ӱ̀@���sq��|�N�m}��^�mI ���.�i
�]�B3��Ԝ)�d�	be�tz�i{׾4e��Z)�:��q>��g"|
���/o�K"�ܙ �'�����Rљ��RU���u�ڋ�/ >�B4��Ľo�(��I�[�9���7��b����C�D��0�#7����"�vz1qAs��g�� ���JI�$�٘p3�ׯ�x��(f�=��rJ��WC�[�MR��*ݑ��<Ck.�N~���g����C�ݭC���M���)�jT��ut[,�<�jR�A�b,J�P3�'���(�	�Wpm_>T
�\��-�	g� m�����<p�g��B���!7qhj$@�g!Y'�A�����n"�R�>~���a������]�v-{�.���-K�	Z����3��'6sO��[�hk�8�1�L�D�U��>Թg]�*;?���?f��0��N��^�@]c-�J���^ɔ ��D �m�0#U���y1��q�Qޅk�륶/Fj��Z��Ŭ.D����>f���u�2z��(�e[i>���� �L*����?h��?�c��	��5+C3�����#`�.�Z�:��1?2aۢ��]nئ�h[^����|
ΘX�ɉ&q_<8E�hM�z����[)mA��y�F�#��e�RlWg�=��Q=*f'�o�� k�nXU�]iPrf����Io1+^�K#��2���u�aO��o�އ��. 5�x^M�}g?�y@d�a���/ލ��2�� �0=�9w���M�ۧ�z����d�C��Q�`4Ŭȳ�M"�/�/�XZ"҅�1��au*��`N0Q����AG%�*T 7��(��e��T��Z�~!�E�,�Y*i�����n_��F���=Q��7�z>?Ê|�#�8k����S�q�E�����4�y�ݠ�saiD��\2���_�Y��kDʢI9q����Wi}+�	{.5<���]v���||�f�\�-��?�Y+�C��c_E�cx�X�E�%�;��3�j�)�g�-�|��Bӥ�)�ñDb��SJ��yI]�T������_[��M�B�41d4%�o�J eK36�K��)�ML�)!�X��*گ���q�#w�"�����`��������5���ф!c+�o&�����<I�1��:�n�Q�6�M���hxú������ot�*Z�$�����z�Q�y��7���0�+��	���Q����orS�?��+˄rǩ$j�R���hX,�vG�=;x��
2��jn�K�/���jYb�wY��y��i�n#�v�!8���Z��C7�Q�f|�������&�*Ѳ�v���Nj���G<�*U��']&������[��"��W��ٮ۹����9�v�Zç����9��V�ƫ���؁z�s)���6��@�]#UM(Gw�C��f:�*n��v�s�� B���r�qs�������~P�8%��P�9�P�0���6�^�xj� �e$�nC^���$���(�8�/��-R5�6xY�{�aJ���/^$��jO$��[ �\�j���'�����n�}�GV���-�	�΅ыB�!����@�&>�b�����nh��J8mG��f�}.�#1��%��i�����G�<��CB)�ʌh�Pp��J��6��-�W=?���Z����q-�g&. ��Z��������FK�og�;�}B�
�j!$��>!���@nϒ����0��ң��UT�j�M�-��������#�	��\XOxa�_G���A�B���\{Ndv�p�����,�T_���	 ��_S��'nk��ût`F6����6|�@��̫^����	1.љ�n���Hci�"��lEցt���d��_h)��qu�lhV֘Xu\��\���X>w�-T}�;2a���3PG�7F]�~�| �V#�["@�@%3O�x��x����)e3�S
@�d��X��[" �X>�V��Jd�K.&[���eQۋ;|D���*���vI����T������AV-�ҫF�U\(*a�|8�f@٬��>y��ǖ1#
YP�(lB8��%P�=;��K岙$�q �k0@�n's��/�*����F"'bL��A��t�ʿ�O�6?ER��s�g���<��v�g��ա^y�n���$����|� n\�Υ�S	�"ӓIy�>��`j��0X�fvXTKy��Y};Mug8\�OI�u�x��D/�J�{7�aӜ�.*q:ikM����xaÐVi�}����I��JAZ��SϷɊ��6��E��,�
�����]zNN�k��|���1���7����V��KA&�_�n���9^z-`o��k�lj�
�O)}���G��z+5�I��g~��m�Ƴ28���+��ic$�@4����.'38ca�-�3��$����Y=�zU�L|�k�UN!��)�A&�0����K���(��B��X���� <d�5�n�!�m��c�"�fgP\��0g-�BFsԝk�n��2�|�� X�e��R[�ӯb�l�FM"����0*%o�nG�� ���l#B�y3����i�2�Q	I�G�B	�t	QҰ\��,��
���!$��Χ�щc��]Z�����H�?��τ\��D(��b��l*
p(W@��w�C�o�������Կ��O��]�@�h���Рc�mcR>�򎗨���{`�]��70$� k��Px�_�n.e]Be��������W� n�Q�;)c���ß��%��q�*���z��]㛬'(�J�pw}�)�<'ջl	�E����C8���j's�>D�K�D���`�5����uy�d����F�G�Z�����HfM͙���X[t��?�+HD��u�0�[�ȓ��+��R��63h\B�)Yt�I��T�t��z�-��x�̐:X���g�O4��z�{�ė��9)�)�Ȍ�݅���ͺ,B_��-=� �!�	��!����f�ߊq�a,�,$�	0u\��k��Z_}}?~�|a�aeYN��v�[j���=�!yI����Ǚ�ᖕ̄ѿ��lL������7����Q½0$_f�@�!��yF����K�=	�O0_��.����Ů
Q���H��{%v�Qc�yٟ��Ɠ�_�ٕ	�5��z 7�<�*x�������MfjG0�k�y��o�E�ʁ��?H�b �R��6��K��:A��y��a������0�?�@�8��D�+��sPx�.���p9U>}}>@�IϧvD��C�Pp����H}皙�1�p�B���_�����iPv�ڶln��X��g<=��l��;�:���,�  �x�U�\/fB��l�lv��N#�A��sf��;�T2��>�����a� pJw���"={��:3�����G��Z�Yx�}ez�a�@F��L]L�z5��f0�R��*ҏ$�O��$�7�\��y���ݱ&$�+0�ٵ4���"W��s���PQ��^��#�-Ito���l���o��[�$��ú���\=��p����{\��u?���VO&|�}Q����e�t4��ѻmM*��;�-�����ND��(�S5	�h�i�}j����O����I;3�1,#W����4�lWM;?��F%RL�N��Ɨ
�phk�����c2E�bb�"h��bS
Dwe���L��@��{B�$���٤~��[���PL~A`��K�C�Va��M<�˗Y�ۧ�w4�U�
�݇��+`��q����빆��E�iuN�Z=_��-�u1�-�r����q|�^3N/����)����bJß�Hj]��f��_���6����u"R�������~6�Z�F`�b�^�v/K�lZ��hK������=t������6�E�f:���nl$^�Y�&6o��c�m
s�%�Z�}��r�ucrY�Od�5�r+N:Bҍ����y��<�^�-,@�������� ��  �5/����,X��o�Tt�[���1A]�fQmJ�v�4����g�U���P�{��Mn~|���<��0�4iB��=���z���
E�~�@B��䭑�T9բ�7�H�V���\�lIHh�����<迂Gs�:���6
xT�����G���_� ��r	�N,�SF��^%)I�Nu/	n`.��v����3�p���Nqr�8�?�фO?�
�"�0�����g�({�?�]�`�Ʉ��Os�+����;Z�z�4���ʘ���]@(������Jv�(�R��_��T����	ǂ��Τx��f�W�>mWM�%�>_]�C�/�ȐD�b�=K߬-6��z�b!�J�4��`���Nc�x����I��L��I��w�����L�7�|d�a�y�H�C14�ÃO��NX֒G��H��6�1 }B�Ղ�7�y#���W|އF�x��)�i~k�����d��|TQ�.���>�GD���/��Cq�������tD^W|-Dk"'�Ҷ%\A��]ɗ��h�@)Q.�&��&��>KQ��v}98�;)αo�9ӡܽī��T,1v��հ�'i(޶��\�򢦡	��65G��-�r�.�l��t�iǫ0�5�z�͐\�0)��<{<r��{�E(���aM4�R�3=e~seA���;��-׳\j����f��.���ʓWx��q��}VU��t"y�h�`���jġ{J2�X��Y��dnz�����Q��Q�j����G#r�j��7�1���s�\��O��2���)�����(�P'��^�^{�0X_g�����+sK����݇�߶ĥL;yۼ��5�G,Q�I ��|���������ϐ�4)��<C��g�Hd�w���p��Ym]!_K,��D�@�P�L�0��A�Z�	$1����E(�Bp�챂�dӻn�#��j�����M�d�Y��Pr��XCּ��:rp����y`�Vz%�g �3}Q�m&�t�3j�-~�hj�4]���9q�HN]ý�k��F��~ح�s�صrj�s�lȯXS�D�z�(Y��y�.��MF}sv;�aV����2d�CR��HDF������dF�l�^5EP)�F_4P=b_�V�h��U6]�e}�~������5KWؾ��3����@�"$������k~L���sQ��-ފ�z@`�Y���E�wt/Z���m��=�H�e�� ��>ߡ�i�1Z�3\�1 ��m�� �hU}�F7�+~It'&�������HI�k��p�Z��m%�ź�1G=�K�X�ל�Vfh��� �xF�ФS����s%�G�@�'�jr!?�MC0�ժܒ2őo��pï���Z���=�OL?;e���yQ4c�SF�[��Lj��QQX\��z��Ɓ%aDEq2UN��~+�+ŕ?Q���r��4s3���1�Z�X�����@]��F���)ͨ�I+*�a�����'��C�K�Š�7{@��,�[ms'��#�K��*�r�6U�n���*6I��n��ؤ��rj�Y���5_�ҧ� H��o{R���{2 Cs�j�V��a��j����'2,}q<��4�4e#[K����>8Y�$�m��'�M����X$C�Y���"��.��9���J�����v��.wh��3�4+g��v�"��p�0�VΞ�����S�2��}� ��������F�:,uw2>���(h�U��W� ���f8����x �J'�z��G �>�N��n+A�"	A�H5��$��w����7���1��8��4�  �`��nG��5hA��wk�,�)��e��Y���CM0bڨ���4�	 f�0�5���,Y�?Y�0*[g6��(Z���6�mō��J+�o�Q}ɯ#"w<䁭:,�K5�9!`�x[��"�RA��������L ��5�T���oi�e�v��*:'����Dv�f����<��%� ��W"�e^�:^���n�����)�,���XR�[�F���:v���v[���ݲ��{lؤ��Q��8���� r|v	�՟�-�;y�x�����Y���Tk��W�iR�`0l�@�r�F.q焖�\�f����i��W\쭧�e5<�2H>�D�"�8��ƣ�ͬ��x0N�D�>r~�6¥�Z�	�vn�IY:�4��3K�`�A��u�8Q���J>z�f��W�B���C����~,ه��r&񚪉�@� 2,��Н��-vdZ
S���V6���	��~�v��8C��w��@��}��,J�QI�\G��Lm1�H�cI�& �7�W��f���U�H��84�-��|;�r
FI��7�P,�Iӡ�ta6��o4�D�u��섋�yQd��<����9�z�=���r{ǀ3g�ħ"�k]��H,� ��m������� ��q\[��j���������;�f]�<ߣw��-���O��j*�Ws�jՒlN��4�.��t�`*
1�庄=�vF����C��)^l�n�t}���,2F��Y6΅����=�gc�0��V�u_y1�1��5JcP�U�Cv�Oq8���3-H���B��5R �eD��b�X�b���С�P���+g!Rb���O2������0�����p��1�l.]� ����CAs[����F�nLh��/Fr��긔�����]��Q�vm�)t�����?�t�r���N��]��zڒ��&2��8d�R}X$a�ã���s���D0N]g��,�֞��|�_Pœ�*�8o#*�(���N{]�q��Yp�f �N_�R=��B[���q4"u&��G�:��e9�˼�}Դ�6�:�9��Z^���.����$s�F�l?SB���Y&t,�lD8"���`��>1�������Qa�Lz۫Ō�6�|pɾ UԩzdQam���5m�$�m�?� �]�i���{.}�&q/�Ɉ�AU,�=<�oZ��s$�=�K�M����/���ԔV��dǧ"�����j��z���s�E.o�
�D�c<T��ū��q�(8�u��n/J[a�����U\۹ѱvvN���#�����q������5] o�����]���d
,Z�p'��D:V�jK�/[��1���� ȅ����P����+P�Hip�n���b�Q)��`ҊJ��H'A}KN�騺;�v-n�����F�4ϼ͐)�%F|r��K�F6b^�Pf�ja�t6����U�ӆ��#I�7S�g�'���䴐]g�nCG�����l���P�+��Z5����S%��$�T([���m���~�?����x��m��E�;m��h�<��U4�gl��6�h�n�Y@뎼�y��r�M!T���9���
��cV�O>�P�g���om@������	���@������7��m�{і�+4��I���p�?;|Ӌ!Ukp�Bsdԧ~>+9��Z�Ct�Y���d�\c�,�����jȁ5;�/�*ct�u��h�5�\�?a���cF4Ԝ�^1�s{�+I�p[�(�"��f'q��[�l��z٘�)T��^��֍<�^1u�(Y�M��56<�׭Њ�N��H��^�m�s@\���1�=Ä�õ��=ۈ���
�}����MPW$8!{�{G�q��랍U1m~Mub��u��]9�*l�5�E��n�.];���1��g�O �TϿ�p�K�<�(��}���^�	�z�� С1��&��7�QF-Dh>�d��r�6ʞՓ5��R�"J������֍a�?I�������}�p�&�y�Vz?0��z��⫊u���EB;3��ѵ��*���%!�� �{I�,�S��҆ ��#���`܎� �|����v����-B�𿥔���y!����_�j<��P�6�h��!P�J{�?.ؿg*<w��M�_�.�6Q��{��2�W$z�|Bݩ<��g=�該U��XV`qW��>�EF��k|��M
G8*JQ�W��T��M�5vU��韖I:�]��X^���訬���{)����^�3O�SX�'�:�C�z]]c�1�]ݕ#`ϡS���`��{;����S=������׹y��XV��ے,*W��9��qp���U�>�':1���?�R�(Ò���|��&:u/_ݙ�		��XR���R�}P���u�c�L\��\%XBH�\>-7 x_P��P�f8狞��r�#Ř����U�LG"�d��S󀞞M��_R�eF�e��d)Ů/A�����w��`���]�����&��=�E��`�����1�^\q莺�f㰎�2�JRL�Y�_�gG���9J{tW��X���8��G�=�D�� V<H[�^S���{��x�9k�P����S�L#p���CC�G,�6���M�3?�6��,����ɨ"��1��gލRW��AПZ���O���`�`<>��Д+��Br�a�.�*�ㆁ�Y|��\�u��)�7���匙��-j����P;�������2į����~��/	���t�QV?5��#j����;�&n� \O��85s4_��(]����D'�n
��N��6
��u�Q��;"u�=Uء�Ŗ��	�U����S��HY���Y�3�@��J�~��/����TF��͒K���yA����rP��)հ����8ʹ޿�@�|
C&���m O+�+��F�vmo
8"q'\�뵑=?��.�
Z���/�yZ��c�r��{~z����?(�M��P8;�r���'���C��)dV�9�r�h%f� eD��
w.P�`�g��p��ç��̷ڒ6����f=���W��9ت������=��m��]�T���/�QC�^������c���Q�*I1�� �%s���B4����.�z�������+saČd�[��q5x*�������_<����~��2�J`L`J���j��h����{����5J��^\t~�ݔ.">���}Q]��SR��&٫���F�מܾǏ�ó.{x�+4�r	n3�/:�d�݁������g۸�~�Me�A��S.�����|�sl��0�[�t���=��O��R9��!0�1����n�ړ�D}ɏJ�|Wu%J�!�����5DnR��،�C���5if�����7-��+<,mb���C/W0��ˬ������z�Fe�;�$.�����`��]�|��+�����.8n�4���� ʙ~p��9O���
��Lc�x���p8>�@��ɄE��7�p�X�z�
���E����H9[�:��M���an��.�D3�5�'�1~�ٻU��3�tb��^܅���P�*5���^��|�����"x����é�B����r�]=��w"�¾#좬d*�`O� ��t��ՃWg}r���%AkfB�iګ[��#�
�֡�s]��ׅZ��=�� ���\F�:'���c�n��AW�#��������Y\CT&ʐm9�ID#<	�d��"�1���7�D�D�(C><7:�4��N;\.�Z �P�ԑߦ���L�ژ	6`~E��aש�NW��/p#S3в*���R�ak��y�_U7�	uк��W1\��nO��Wz6�{���r�@�uNB�ɺ� �x�+��э]!1�'�s�1E�*�It0́:��Z���/w{����΋�¡Q���Z,Q�]t��Pb��-�)h�v�l���l����h�	ڏSx��.G�W�+���b_P���3acC���r�"T��L����+�GX��~J�����`��_&�]�an=)�m����� ��>��]^��F�ŖKAh���z�

w,*��[ ���J��:��t�D�$V���yG�2P)��ݱ�� ��Kb�=_`�<X�H�l�M�G��ܽ�EPKO�8a��`�����V�T���u��Z�M�^���"_$��{�#�"�:���ڊ���g���u\"j��s���������8B��[N�N ]��fjbѸć�btf{FMb9��g���5k�Ť�@}%N2�֎�}��b6���O������,�U2Q
���x�g�aѴ�,![�v��ܡ?Q�Y/f/ZPf�l���Y��fЌ,תqhc��)�p����U�B��0���&!� ��������
�<i#�M&c���
ϵs�FG�d��1t��y��T�����/�|��rn0%6\�/V���WD�}&1ˍm��r�u/uJ�`�a\X�:�t�X�~%@�tT����%���>��l�)��b	B�&y׀�$���g��-X�9�jAs��'V�+�i#bL}��.K�F���'�4:�ʋɚ%�5�B�r�Zة�w>c�̊�|`����e�)IR�*c��ʜw��W�{�z�����gG���G:�I�)t�Șc��͡��k�˖�������dl��Ɇ��H5�3��3x�U��EFW�Qb�ɌU����l���(�fS�=�2�3S3&��Z��ʿE��[��l�}R��^'��� Z`�s�dq�pe�͇��c0=[yqBn�z��I���X�^~M�og�	^�~�3�)�Έs�����e�#sߥ����D�پ��nrI��+^}@�us!H��H���<��  �����Ae��P�!0ۊ��a������]�ܾ*��YJ-�+_<���(�)Z����n��oE�ҷ��'����q�Yc':YrktwD$��Pzw۫J2�͒��Տ8c}
~�L5��1-�9^u[�^����}�Vgò�Q��7M�iP���K����t�,@sV3����7���,طd����A�*�+g<�$�F�s���^w���Q�?Q<�Zn��Sa����%G���}�\wn�i@�[jj@+��`�h����0��"�L$�t�t�|z���0�Q����y���F��_�vc�4�%%V ��P[)o.b�9�l63{U`�~(�����=(�s1�O�ڎ��+�%�Z���p˜_�ѷ�R�+��\�<�������C�Ϙf�R�a!jW���#��8j;	 ݯ�\uӠaL?��PC�8���f+9[p��(���7�XcU!�
?d�7�2^���ҡC���y���%���ߛ��_L @��E�|���\{ɍ1�����ƼZ�S�[N��������[�Lo�p)D���6�ϔ�9<��'�t�~��\��k���,�J��Z�������N���s����G� �a]`.uo���jհ�ų3�M���o-����t�b�;����
��u�焵he�Ǿ).�����ʤ�slIk�m��19o�b�W�d�E�6�^:�pU��2��Y���&�Nu�}�>��<J}��{&�+U�����mz [	S0�Ee�zh��G�]]��W ���W��gt��M���j�A��v?:�%�E�D��зK07�$ �h����VIY�xð�<@�$,Ë��d�<x�uu�k���5 =Ϫ���*���*�l�����}+*�_4�|���ȂŌ��Q�pc]��cӗy�g����:��Aj�-�h�Lq�e@ϸ�/�L��Hk'�W�?�����H�������ݱ�S��.�����2�؏����1;����t"2�_�����ޒ��U9��x��wY��V(����J(����=��� �k��-�y�Ct{�sE�w��2i!��0LEf^Q�2��5��ʗ4lm�Mt�9T��}sU4�<�t$9�W�<�	Y��;3��$P��҄�^xТ|�ֹxZ��ES�_JQ�#�K^<\Wca�`�cz��,S���;�����~2�@j�r�!Q������Q�s��Έ�!!.���(�8���i�X!�P���6Ћ�>L�Z����Q;K���Bb����d{���Y��3�c�ut'� uG���ڼK=�ܸ_�i��H�nO�8!�����9_�egO{IR��"��#ȮX�����}������A�b_3S-�G�0�,�d?�n-K}[�nQ����90�p��#�ڝ2?Ll-I� ��`lw�
��)�xa�F�!� �«�"�}s7���X4M�w[�n� �a߅�4Q�w@:ĩ��F=A�vp���_�9��\��3�\�����*Vt���CS5���������?�?�&���#�>��+uj����Zְ�=�HV�w���H�zК�V:���&�C�'�tu]Xc(3 S��)�w������:��*
�W8#WS��"e�����sg5�Q�������K����~yO���W�Px$XH������	�M�ts�)�K���g��fu�	ɸ�\�Ak!b��Wnk�s�h���OW%�lLL��o�	1wOd�������J4+W��:j��ɽ7�$���2��B=Jƅ��3�&�l�#_F'�IEw)�����s�٤�ϫ�q�֌Ӝ(���59]���\)J��zUh�6R�{��{	����`;͖B�~�ӛ�S��v0��6�3��
i�\�`���2N��s޺w�϶=�(^�KY]e�`h:x8��D������KnU��=R���YIG�&�'u�s�lL��x*$�=k�7��V2q�{��^����ʂJZ�X��bW���)�[y-��1�屘` B|�7���ȸn�>ӄ��`�x��u%��u�����>ù��gR9	��a�q`�����<����i�:��k�n�;�ک�6��A�_�UUZ�C�P�7} �8�emص2��L�o"�&����-�W�8,��];�dZFIfiâ���8F�B�`C�U�8��P��El[�Eo��OJP����c�|�2�s� ��	���'�7
�e�(T}�5!{��k�$�$#ȥ5Vy3u�����\�\��.4G<�=D���n=z�j�R�����~{b��ݲ��=35R%��u�������K�^p�9<����m��5��,Cb.���\s Ҏ�:*���U��t>x��
0���l���?u�v�ղ[��N'W�N�S|i	���,�Tl:5���}`�aĥ�/�j��?��;�P{�I�j���g���;��
�h�>ڵ"HِK-wH }�C�fYi@)�ߕ޲}���[{]��.mL$ˤ�P�9PN�#'����zσƾ�=�͹'��CKy�PZ�(6�h��)).#~M,�֗�&ڛj�)d����i�+~)�l�i�%��f���=���ͧ!�ݵ�L��	X
_.��~yx���!��^Z�X%K6YۘӾ/������o�ܘ>���<�~N��������c���Yb���}+[ V��ոG7�<�
�}����`��Dc�.�}k��Kuoz7nj�n|e����&�0�l��M�#�A�V�f(��3�[O�W���a7dǻ�P�W9}�=�]���O����zb7E�lc����'e���o�:����-��@"j� �o�x�O�����+��P��&�����Db+�>xe��"�'rr��&!0��_���͙�ۃ�'_�c��%b�Q�\�c2R�14�ȅ�>�3�F�]���m��S�:���<���Y�˃�7�<�M��J1]"��]7��<Ȋ�K�� 
�R�l�H$��)<�@�����S���I�F+�Qڍ�� �3%�ܧ��n�8�����
mʸX�"�j���B,��q�!���ϡhQN߉�fd��y��G�~�'�D;��(���&� ,QH���FQy��4��-�����������X�����|E�包0�hyY�,t�{�u�/�ÈbT$A�u�u�\�rh�K����VL[Ab��(ױ���3��&��[h��u��+�=�=���ͪ�Xƿ}94��s���(?�k�8ϙ�׏���0�w��7m�J���o�"��D�ڊfW��7���2�-Lu�t�g�b
.ѿ~L�n bl����+C�k�'K�4.�c���v�~2ź���d�Y/��-����?�ـ:#��t���P����8	 n�A_P��2�� ��fߧTdəl��2�R������ح�h�Ԋ�K��3(�e��P<�!���V��|�!C!Eb"��]{���#�>9ô�V������X#� ��\U4v߅��YC͈�g���"��� k�E�V�@ސ{t�s�*`(o�ҁ�T��P��[�Q���p�k���|��:c���"/'���NԓͻNח��e�Z���@	�*��	s	�+�:W2��@�4_��}�ˤ����k�����FCB����L�ʏEK����$���v��K�*�T���0�Ӯ9:�CGl��+V�c,e7�by��g+D�D�}Û2��f��C���&YiŴ���o�2>�zl-�
:��`�������� �8'G7}�x����bFA`\
�MX3#8������L<TDS'��.4�I���+���2Z�3�D&`}�-G�Ă��G+8Q��s�;�G/�8ڊ;�M�yԡ释e;���~�&@*�mW]�ҀE)�']�@�����Ŏ1!���H����$�1꽺�w��E%K�����6�� WN	PY������ �r��Zꈙ��F[Y)�%�^S�B�g��&R�t�θP"晫���|4���ғ�[��S�V�9!��������F�rK�^Ã9B*�B�I��w,���0���P8��͔mE2������y6�U����2?�p�~ј뫎�Z�� VE~�0ƂQ#���C$l5�Ř�2�)�
��A�s�w����J�gA͍KST��Ok��t�x�0؜�Y������t�Q�<aXX�����n�R�Xa����3�V����r�1a��&UDxv*��j�[J���F�Z����!�	�nb&&�ܭϊS"�G����K�����`aCh�(Em.���p�dJľ�I(G�H���_�.�6��!��C(�P%f׊������$qmՉ1���i���{����Ů�L���\W�vD��e�+��$骫�7�-܏�G�Y,QU߅� F9L��v]1k�R���ja`^[6�I,,:[g�P�t��j-;�4;K2�[ - "[_�Nʲ)�BIY�4��a|'�Ձ���4�6I��NXZ�pA��g�O�>7blZ��q ���>�.<J�¯K{>��9�k=��U���7~�%�E��}����Rtx>?���e��eYRѭ�RߑƉg>B�gB��yȝyO)�䓳����;̈́���\0K����5����͌8�|��X�K���9Q`�~������8��*���v�r53� �A�x}'LLQ��~�`�s],����!������5�X�ݼ�MA],��p����G �Z7�H�p�M�e�d�[��k�����r��b�$n�!l�"]�j�FCE�OzMZ0����Q[ZRg�_�L���H�Ue����U|"����vQ����s���ݩ��]��CF�!��6%j^��A�Tڕ�.���SZ����X
-����
��A�ӱk*�J�=x��ͷ�J�|U=��p!��d�)�͸�D���¢��BTM6ƈsxq3���El7_=���aj��V��Z���E'k�Ʌ�Z�� Y1$���]��t�T:�$��ʹ��ў`�~�K��ʹ�� xBO1����0���e\���5%K�ч��_9b����������D��$ې%��K*
�f�#�ɂ$^ϵ�F��f�Bc��	ة�Wt�f�/�n���y�;�z�aH�����""�os���ƪ�iL�@��e�ߖ� �u�W�i[D�M�u��c�4FH�:�����1a�R�F�2
��5�6��x�n�����,��q�!��hUC�~-��6;cPrۮ�JA������\�Ռ�ҽ�Q��n*�$�r&�S�j��H6�;��~6���(Er\U�Kc(�
'n�����q��I�ޣt'����y�=�p�\��MR��>��+wi��}����%���<S���9_V@HU\ W�ծ�|�%jgV��wإ�U�=��U�}Pݠ�:P�z*6|04	Ƿ{�� }4E p��HN���|��ɡ���e�w9~����J�|�;��إkZP8��	��AE�u1�n�����B}�Ga�P�}Y$���6,�x��Bxj�N[��I͔^�Z����次J>�KW��m�`@.�3q	$��[CC�1�,���;.貂�N����5�,	�'n��A������>��M�֞��a������/��T���s9O���0a��;�:�hn�ĩ�L�z�Et�E`���ٌ}���hR� ĺ:z9IC1���ފ��PbaS_�+�}����T?�����&]Fv�"�e̠'��Pj�+���@��,�Z^����B M��Jm^ʨ�x��~sm��G#"cw�d;ڤ��q�� f�!����)��� 	���&,�Yݓ	����`T&ќ�a喯�,�rm�4u~+��S/��]�n�
n�յ7(x��C����nXd��;��3�D��Kv\
qȇ3I[aB����s_�.m��UD!�<�{%e��+�K��<�c6�2��I��n�D�f?n��H�n�]�&�iVc����B���7[:��1�'�aO)�6�@���t;ޗO�s"	tJ��)�v�o��IȮ�G��x]�^�G�Q�v���U�ý���`��Ұި���'����/��Yo�z0�Ua�+t|��ӛ=c;G�Q�sxn�{9<!�?\*u�,U��kD�#��GI'��L�E�,��L
d �������;m��G�n��*��%���m��H�.������P ��5��G$.)�.�޵��y�|�"�>�K�2ù�����*V��������6$��o�4��U�|UP�0��爤-Y4��$�i�y
P7�h�eC&�6���X�w':EC�5�e�_v� �М�+�p,��zSc����D�(��a,�ˁ7����P�P����z6����{l��.7]hw��E��f����t�hn,��d.�X�-�0gɄ�+ߊ���`��!�����9�*��C%˕2���`�Yեӫ.�� � ��a��1N�r�M���uV�+8:�U���/����%� �������!��"^Q1��d�1	�
$�L3��+�d��\Z}�ߧ�9�>��f[l��6���gE*���,��ޏ>�h�\�o{O�3��9�6��'�}�)SB�;���&����.!�Gl�J���{'������#�@�$?��V���®m<4{�O��#�<r�b��k�X�cƦ���#abd�yz�T�����|��g��:����������f&p5�)<�C�E�c=�~=v�Y�r��@��zgex²O�,�����`%��o��*�����v���s
�H����N�0P��.����Y��Rw�v�����!SJ֪3��}�П�����m���l��`j:_\K�E&-�+�n�B�a�A�&V3&��	�ʦ�����U�}P.49v �O���a���EZH���&q���ؤpX4���!���-��W��h�&����b�V2&��~�:��%v�)�l��_H�x�޳�Օ��z�o�f��aw:?�n��ũ�r�><L�ED���"i��D�6T�_9xR�;ŗgj��0C\�I�P�|�P�L����/�,����o�ߪI�ǻf��y�e��f0��X���dsn�%�u��D#�z�+|a'�E�d%t�2GU9K�x1�<RA慨��g$5����u#�b���!T�߭��|�M����ۈ�*Ɵ�Fcb/6S�S#|9~�չ`-�,@=��
!���H����CC�@8N�����⏎���������s���b��RQh�u�]�(0u���i?3�7[x�A�d���C�9v��vcu�]�^g#�~�5�� �[�h�C�2}���ԛb�%�j>:K���a��EO�5�G[��L �a"qK�y����<dQ
#�������<�?��T�W�Sz#liY�ڗ9k��g�}��rl��5O�<� �N�y�:�����_�G&׶��P�W����K�!�ա�G_�W�x�"	���RZ�ܾ����,ΏI�:�FTw�b�8k!O�ζ��3<Ύ�F<�x���[��É�k��9,��̨Y��`��]�m��O�:��<ʮ��Q�7ިl�b��������6�_��v�A0!$q<1p�0�U{.�#*�id�L��u�|���O[��@1�JH��Ŧ-%vwB���0̽�3�����ԍ��?_%@p&S��;k�L�8��*��*M����~�
��M�$����,PH! �S=�#Wb��$=�
��Q̅�U]w��A�.t.N�׮a��I2�끴縆�B�D��K�R�G�`l�* �V���I�Z�����ZI�}���ow���g�lN�i��n�-v���1��?�ba���g�N�j��ܢc����>���F�bW>=zJ����ˊ/��Pc�D�j�Dd
����R�}șs����5K+�e|D�� ���I%��%��b��>���i�ny������Į���+�`�J�o�a����ܿ#��	��oU��Ѱ^F�Zg$���V��[vM�\�k���pl�,�9�(T}Yy$4h@��h��-�v������!�/�@w
!���^����l)�<7{7���\)7��\n� �m��`�"]8u����P��z4k���Tx��"ɺJ�7O�W�68}k�p�s���q�M�%�ܹ.�4+�d465���h��O@�cO�їC6�Ȇ��)J]�f�_2|�����dI�ɏwI���M߷2o'��ά�>�i$�]Fz��f�G3mg��K���ТL.��AuD$�d[U��EҾ�p�EP��Ɓ��i�F&�]���X%���'9���rx���kk���u�����Z��҄��-z/�ܰ�����L-����$_d��	=�������!kF��~<�,�;���U�gSFi�B^BTJY/Zۧ�J��ܓ l<���hx������l�nX�M�&E
�5�#� >ޢ(*�ϞY���C�r��`08���jks�Sx� �Ěg�a�Q`�k�hmAI���A*J���L�T1���}"��3�R��I�-,�b,�Z�Į//�ʮ���O�0G@d&zD`V�"(L�<��c�,�� ��B�M����ĂO�wאt��F��Ծ#��}�jF�E�ۚe�B?X�Ε��v�_���!o64�`hŝX�s΀�/2E(y1���{ҩ�T?����X��sybF\<�J���䚒Vik$�v7���3���,�hX�b�º���#22Y˔8�]�u� �_����g�7�|�i;<�q�R
�ɓ-8{��u?���ØZ���RT�6���P��U�BQ�6�����rq�8��n�(�Ҁ�Pav ���ԉ�bT��M��G�j���z6�2Ђ���U!,J�[4���J��1�v���ez�̤��輕��(88���,�a�ص�N�����?,�-��)���]~m؀��H ?�aiB����(q�Q�E�]�K��؅�-K'8�,���[�k��������<��wWk��Y�����/j�U�Q$���T |<EK�i���a1���I��j�	��<�����PM�p�ÀYO9�6��>2������HA`q��L}��A��r�ʰP��Ufh-=�g�h��PG':�5(����)�h�NT~#�������cK̀��Ħ8���؆�������ǯ�<!Z��f����*v�F���W�|��D5��RK�Vu����?����[�Ms�4�@=>�C��"�;�fIow�]2���a���i�t�W�'w�����bs��돏Fŝ�Gn�ԧA�6�C1������s	/fċM�	�-9oR�X`S3���N��~��R^�0�\�u�7k������Ll���:��{���|U���nP���,�AZ��dEk�҉�s�a�u�{s��?$�I#�n��X3���1<_>i��R����Y�����adzcA��#�vy��� ��V�:��w�����z�}=�w�y���<�#�� X�p�����[ʪ��h�z�!|����1��#��ޛ�.�1�*��y�@����/�X`�Z�	���7�Z/^:�����%�����"j�Nr�~S����N=���1!5����Jxř��ꜞ��*R���ٍ��ߌ�9�>����n7�J�� y��/S�N��Q5�����x-O!�S�)��9j��L+bW�QY2�8��^�(�S�v&�ɓ$rq�7ހ�)� �����������`Fu%e;�t��ᬯe�.b[�l� �Y]+N�Q��tc�$���g�9j�7�cý���S
؆9j���('v�>�{,��HZa`�A	�7�4�G�k%Hb�&"b��K�B���.?��	ʡCx�9$���)�U��Y��;��*�~ ��.�hS^N��8�Zr�⽝B�{:�m�M���B>�'Z��׎����ܘ�~��>-�.Nm�H)�*~L�I����~�0�
�{HD�yx������J�"7@�0g��W4)�[
��Ʒ�د������ �a �:5[�*��43�%�l3�E��sq2�u��@B���{�B��{/8V2������	ayw��}T�DS{=�=ޙգ-r}c�Mw�}�Q����r~2U��w��/�YN�Ϻ�{��?��q}�p/�WE$���ů��#��5�mf�R��w>�#��J�(2Q�~����j�ŷ����6my��*�$p�6kb~<9�i��J��/�2��b�z�Px��iB��Bp��sߔ[S�������l����(;U�W�YG*��>�O��v ?΅d��o���9�'k8V�������TO�����wXBx�?v�`:U�4
S}��§l��{'�+�w�/���r7�4�.	�Q�6C���:K"@��S���Ά������!$�!6��ڥ��
��<��=��� op��E�P7����;�7��=����RŴ�js��P5;5�h���y這�LEh�r�#r@�|Mu��C9��2y�Y�*%?	B&C�
Zۧ���D���Z��D�a6�<�!j���|Q�t3-X�~@�8D%ז�e�4��wjr'w*:��nO�����U�`;k�������T����j��-�ֵ�����⵼�N܍�q�.n�B���8sg�iX=#��p�I�T��λ� �ً-����%����G.��b��X����64�ȇ�M�Z��+;d����K�87�b�q�������� v�_
��t3٧��\p[2p� �T�ÃEG�7��{N㜏;N��/���4�H�A�Ĥ#��JF�պ�a��������/!����x_�S*�G�����[&�.�$��q�^���'Q���O����壹�N���g?���7t@���Mv����j?x�}S�6����G�+9�6q:�h�FE����=��M�A�J�J�]���$s��$1�H�'�Kڍ�sʣ���w����	�# ���X��=��� I���{�<q��� ��2���d;O�I��n/B���v�L��U���+�ַC��KɅx0S�)�T,[�.9�������R1��?�;��"qq>�^��˱�}������_oG#b͎��g��<�rr�G&�)�5�w�y}W�o<L*vi*���&��1Z��NK���A�$�</Uqa��gN=��ѩ��N�[[�A�f�^���� ��1��ܘ��:g��� {�W�"�$L�9�d�)"s$�um)I���_�����fD%�z�N�����9�4xČ]��� �5�՞<�q����o��E啸�vU}1S� >���c����� �Ar���/L�G�`v�	1/︲,^��͇��J�>����Xn����BɌ�3A����1��q�B���۠80.��"���ֽ��x�BB$(5�cH����,��e@�u���Ϣ��0�Ѝ>�K1����KBL��Kُ�zk.2�.�=�k�,w;�a.���`i�b[)����8)��x��a�� ���8�u�+qd�
��_�7��n[.�06B� ̒qw��)���;VM��)��ٟ��=��Tv�\�
���$Iϟu>�|���H�=�иg8@U��V͉܃�&\~}��\�Ϝ̯E�|��ޅ��V��^>�L�����֧�M�PۤM��"ϏO�e�ԉ�N�9P�/���z0��2������7}|.\ӑ�\r����Ƿ·���)8�Ű5�b���M�@'xd�*U�Ğ���_�N��	��.>Pg-�.�ٌ���X�T4چ���h���B���d��&4����G��P��z�[��f��J�<v\�@�
i�=��t���`���t����Cl��u�,7�M��Jܮ���T����vJW��ʝSIzީ{-��V־�c�_p_��Lj�F�W�e��X �Bu\w��΋˄�B�sZbJ˕�m9�S����<}��<ˁ�H�0y�bpL���E�/5>D��奏5�{p�;cr�jv8�n(������"�4j8f.D\�� ^�!��^��&��*��_�@.	�1�D���(,�Y��!?/�k�pc3`�" �@�����"a@TA�*��7�[y�#t�'�g�qXu��ST�Yl�W��k� �	D�l&��m4J��.K�[���6yv�<Z(�^᩼T-����U�j������0�@?��`ghjRx�P�G�t�5�gwt�,��hj#��ӫ�i���#���[��|�s"���{O��H��^��U]~�p���&�&��{,*�g��F�ar�����G�O�6L���|�	��[��o���UR�����"���M�!S�-H�	��R�]��g�����q�]�ք6Y]�p� eF���r]�FZ�5pLU�У��+��;�k!�v\����s��0���� f��dt��S1��xC#����i��?�)jB���Vؙˮ���7��Ł2�WM��W���{Yϗ]��O���3���B���L�q� +f��;�V(�h��5��,�3k�M+$z{���,���}�*�g�|��:����V�0\�<����y��C��q�c'CƷ�&e�/m*T[l%4�����	�])'�Øa��ꄜ.>9�>����e!�B�2�\�7�q�t}k���cf)'�B?�mDHX�k1�D�s�i����Ca�\��y�".�tRd��L�-�B]�����	 �C�y(�^��âX�,op��^׈3D_�$M�1�@S^��82����S�V���̓^��!fE@�B�IT�@O3��ga�.�E��2�l���?�Rz�Pu?�� �n�4A���Ȭ���n���>�Y2�ǩq�]��11���7��_X=��T�p���BD����?����u�m����hc\�46��݌(\,��U��`����j$0��?W(k���f{xe`�Ѡv�@6��J;�T\ia�x�B�h�$HT�v8�;���7nH�`	q45B4I�1,� �I������)�~���&�{1����j����R\a�Z�������(3�^��'dM�FxMWw�9Z*Xg�ņɛ���k�5F�fv
�BW���֍�)�`�}�J֣Ϫ*��Ɂ~Y�����6�$j2�>�ر�K��#K�
�أ:�$�-�ci�_���{����p�K=���`�(�M�Y'C��c��w,�zSnoj��7���zjwyn)��"&��d{�`4w��n���CZjdk���"�K�l���R1��?�7 iQ��� Mw�1o�M_�/��P�'�O&��F����	�~H
i��0��Jo�&:��� ԩ�����Js�ܲԞ�ՙ�"�'�t`8�E7Q[hõ��UK���@��߆��$g��)��-���̇��mN�R�j&��1l|��Ow��<x��jw����WJ���0ۀQ����	T9�_��wF6���|;�0��!7���4��˅�ª�N�K�59�,�Q������l��kh��R�����D��
�#��Φ4e��'W�4Z}^74��8ڪ��'����K��E�Ft��l�B��\F��Y� �6p�mc�s�7:���_*a�;L��]�� ��=��Ug�8X�q*�� m�gq����5�J�ZZT2��߄L��P!�HL��35�JߪRp4��l��G�X}�ɘ�5L,
Ԟ�k3�;���7D�ᝬє �Y��ݖ	�$)0U�M/!��[�\�cU[љ��VĪ�@t��]YR�u�S��k�WO}�5�U��x��tx����_�G��5�L�>�>��<?��Z��Eg,��������f8X�����+��w���dWa7kE;�֓�yY������H{H���?�_}���[�x^q� ��%U����
2W*�����H}r�u��
�4���4(�}�c3�ͼ�>.N!�{�/���L|�3+���n���V��l��ˋ��9�vbn�d	@h�1�����<Onp���1}���P�T��|�9-�=�K� Y��L�D%�-�M�е�d�N���8e,?Ė�
����:Ɔ�ڕ���'�tK6 ��bu2u� 5 ���[��4ؖ��V�� c��� :�Fx��b��u����|��d�ʫ�CxA�y�7��Kt
�RG�Ts3��@��i����|뎉%�IX�u�dCh;�]ń�H�7�9������yx�����$���a�`�0(�H�5��X�u2�:B����/�J�ڑ�R髏��������,��KJ��=@��Ե��RaY"���4[�	�[T�F��C�4��z+#L�\�H�Q����;�f���c�~�W/uѥ,�f���*;s9\n5	l.�:x���B�y:�R~B`�,�7i��*f^�O�e�\���kh��(�*f���(�B����b`BSJ2E@��sF<���
���!��R�M����_�~���"
���E�L^�Q9Z�'�J'ıC� �W3�11bhF^�Fa�*����#,͏��O�p��3�/�-�rl0|J����B�;b�me�x��^�,o�>-�?�����������0OC�yX�w4V6D����҇���ُa�GM���]������t�>��x��u���U���GՔ�w�ӃxG�:�A����Z%UO�\�(�V��U�8�[�d�y���F��v�AM�H!��2OIv=oh���$>�s�6�4�A��$ hP+{Ԗ��x��5 ;�0Cu���S��ǵ�.
���k3H�,��X6�/Ew��c&B�#�yc�@c0:�����X�/��-2A�Z,�Χo��ߤC�|��_���A��V
W��� �Y*�c�㶭*Y[�ۉ���D��[ҷ�v��.jLu^�~����ߟ�"�Wv��i��� !�#���g��ӛu׃�*��2��i��L��?��S�清f��NKYσaĘg}C`VW����7��`�@�ɀ�i��vD� ��vXg��-Vzo����W����x+J��b.?����\3Hz�j���!bt2�Z�e��>z�Ah�y�w22ri-*�_�$��5��{"�q�uUW�������<HǠ��s޹�z�j�:���l.�//�'D��L/�UN
̓�J���絓�<E%^�I0^��)�|�Mی\)�"��z����l66d)�#�/P����Z����OX&e��)����B(a�t�_r$��53ҭ���p�{��g}�6=�����5��-���Q�F�`�mLɵ�i78����梫*�4=G��}���d�J$m����[[������HJ;l*�*�0=�&C��D%�k��`�I���꽨[`$Y���A<�S�P��<2֑����Ncծ�^��"�Z,�\�R�:���*�FK|"D�;����aS��η6���hI�`������v!p�ނ�,����j�đ��<Wp{-�� �BN��c�%�֝u(5>s�G[��>o+�JU��C��H��	S24�b��
�͜"�.M3��k�W?����.�;)�,���Ɂ �b+_иbr���[8��w�k-� �D�X�
qߦ�U�*��~��\eNh �]����A�3��p�y$M��nq�.�t�@���k%N1�h����~��c�@?]�xC֩�|��������'Ų�$	R6�nR8�A ۏ �5��ݡ��r4'b@��=�e�S�3���zE�@*��S`����}�c�D�M�{�::|yA�n��2�'�Y�nG����3�)�2��Ɵ�cP�����pوe-yrϛM;���%�d,���0�A&F_�^��2����<�ѕ���@�bhLS�Ǵ^/Z�>f�`�<B���������-S����`�?ɫ�o\�z�k��)evm5u�E�#C~��$*�ynT����Ţ�!��Y�+S��C@)TX�?+|��Y��u�II��l�ı�R)�C��Y2�JR�l��8�1�k�@=��E>'^i���c��KV�H���w+�rwR��0�qԗ��hf9���U8U!���u8�S��(h�"iI�_���eS�e�x���|@��w�)�`1S���X����/ 17�ڿ�F,_?�� ��	З��C�BϹ@ng�[V�z[x���duXMkx��$����r�lP$�����ݡɓ�v�LXE��ҵ��ud���}=K��}EQg��(A�uS�e���b���X+UR����$���	�%�+���)�����'R���Qޖ����r-�@Ԍ�ɑ�[8��2�?i�ԗ��Z�����F5��Y�ˆ��/�Sw���7S�[&�K6��P�tT�h�Ο�H�**�\��4����+Ť���|*x�-5=�u���sO"Tv��$��]��;��.7e�J��W0�,�l�<�9�M�����h��k��+x�1F�w��#+i�CE��Yk�$��D_=lx��',�&j%"J��2���Y��� ��S��Q�����K55,w�t�}�]�C��f9v$H�07߷�ӟ}��tq�2����=R���n��gc5S)3����t?5��z�X��3����xn�H����m�j�P�=p�{�'�@F��؞����z��>L�ϋ�����5'0@ǝ��N�Ĳ#(Q�`����t;���3���ح��h�p��c*�z�� ?�����\рѧ2�8A�7��W���R�T�mǱc�#u<� ��0���&(�S���nC+2��nre������mT8b�K$���*ZP�JT�ܚd�Y��o�ġ't�g�͒(ܩ8|�	�4�=r�@��(u[b����B=	b�SrI^�3� 8U��~��f�
��w ������ocXL	��H�>�}Կ	��zf����[r�̜�+:���t
3�J+G}�����g$����B:y/� *Mэ^d{7�nX�f|���-��2�A�Q�sIYٱniJ�IU�iu55�ˆ�JtdK���ӭ�Q-?��t����B}��؁@�h��\��P���7y���Pbo�f�q#�[��c�d]����1_+WA��W;Q�ݧ
�G�����3�Ț�/��c�(���)��:V�,��������{]@�e%�q��A8ɻ.��b�z��`����R�gf�Gd�\Ә��?5�q�ƞ�ç0s����ˢ�E�'�N����5�D:'������BR7ڌ&`����9Z��y�th=��a1���D�Hb!q�w��)x�^���"#1d*�;n \ƃ�[�@괘�0Q?��qRP6����d����9in��Q&I�*;�����xw7��bG�L��X�b�� B�����*ؔZ�:��[�7�{�:��rzyg"x��@Y�)�d�+-V����l�0��W��y��g!"lQ��<����=��àA��X��T!v�B�2�X�:���q��ڦ�?)����2���;NS�5�ccg	��+m�X��Ʈ	���k8Aw���0���'����X'�lvJ��Ǐ��BB�)D�u���g+FQ�&�Z�&~���$-���}�����8��뚍�O�"�/�f½�/�5aH
��n�|3�n�WmR����D��d���CX���g��Q��<�pS�����8��B~��$�Qt/!5
b3�^u;�4/���p�i�#S��ۅáA��+�2%|��)y�ȏ�Nt~ɢ5��x����2U(�l��+����5,T��"����r��ڂ;m=$t����t�[���6���:��I��_Y7��B4Sk'�f�lj�������`���&/t�����/������m0����g��7ʊ�.����d�&S�_m��s��%#�{G����

3��D�8�8~��k�T1��TJ�wu��u�����>c&���VX�霍@�������j�4y�Y��4�T�lApC/K�{1�ǂ�?���gY�p��2Z��qu���?��j��e��Q-�4��
�0�g�)����C�Y"��-�+C\%���5�bV�V���F��_wCܨ�@g���9�.0.���;��_�/h���s��|=aE\"�	t�b������Ta�#=̈́��`Q��26���������[�'��i�N���^wB�b�B�Kj7��7��H�����(�|�y4�Tc�n���8��\%��o��ȹ��v�>IP=ƕi	>(['�Аd���D�.�,'\�>���mD�^Y�d�H�.����G �jR6L�Z��F���n���u
3C��u���.���X�:��-����`��z�e��O�B�r楌m%��]�����2�E��ĬXrP����a�ku�~�O�IIu�m>�^��7�`�(k�������ѱ�R�1p"�,� {����y5;�L'&�����~$y߾�
�2��6��cw��ze+1.�쿎���-����^Dz<��8����C�X����#t��K�A��,sZD���+��t�:檺��>�7$����T�N��иȥ���Uxg:��MF�� F�a�=��Z����
�4^�
v�����jT��������E�����\}L�uQ͟��F-iZt��׋�����e���	tM{%%#>�a�%����̓��pT����/l��⹽V���d���~U#�\�g"廼5N�D�^UM��0.񝦄���D�#B����uv8߀!��,ۈ'����brȜ<��2c�pxY� �p"p�ƫ��=/��St㹭�R�ۦ��{�l̽�%��^	�����$�"T*����w LW�[4�%�Y>�+����~=Ֆ�����@e;���*���"\z%2Q`�L�Z�1k��3W޽��i1ݱ5�މ���*��b�s�k�/.���p�b��)N�r��R����2
ț���q��J�x`&��w��F�ð��]���k;EM��׽,��Gf�`^���Q���5�d��X�`�w˱A^�ሊsQ�m�|��C���n��Uw�f�2R��m�@#)~�J�g��\�u�8�pj�]�=�͐0�E�Mo7� 
���Ζ�'� )m�>-kn�X�yߕOd��i?�z�Q"=�ʼ�;(@��D���^>j/�<r�B2\؍*5p��=�:�&�|�����5����������"�D3L����l�Oq5@B?���q?�|}�ӇĐ�ɟ�=�C	?q�
|�\ �p-��@݇�ycP��+�i�����%{PIם>��D�O�2����λ`c,%�E��r7���Ը�{S,S� ��JK��,VVk��,5L΢�������*�<�kP��1�W. �]����]2xM��4�O:�o��Y�ذ�V,[�ڀ$i�8\y�y]u�0A�9�K��`��]�D���du␐�vi˹z �ݥl��m#�kgR��RG-�����H��0ƹ�����'�W�x��*��; 2�1�ի��)�n5���=M�R�>r!e?3�iD�NL>��.��6<�;\_K�tb*Z�%J�7��!��9~k�)���Y� ����!��ŭ�q^iV������B��/!GS3�_�o�K�f���?~����Z}#u�}CUl�=�c���ߩ��b�Ȏ�2��W��?�4W4�頃;>���*�\����.�va����b���$5,R��Ͱ�?񯨵JW��nW�x�ߊ޸I�ٷZ�F��r>�b~F7L�w�#=���y�K\�a2۳��Y"qpN�HY?#�S+;�/>���5�O�uw�_�SѨHCR��W�ؼ����s,H��Qo��'��xM�Po�.|a�'�O��fK�v�/z7NGw��z-��lSѯD��΅|鬌x�Zc�(�  x�'�N���Q�>�_a�Dy��D�l=Y𘖥I-|��Ì^����U/���������D�n׾���$c)��~�G2�f�D�֨c�+(l���/�@tI�i<�z�V�t�����(�6G��!�s��`�/p��W���$�S��)�v�r�N;%ĪӅBW��w{����I�U�L.��+��fG���!��g^�^"���,U�!��0Κ����%��ë��+��;��sbg��U� �VE��B��s��<a���]�ww������f��i���6C���@�ߊ�.�q���2.-[�cz������RN8���x�?��9g�	��~ӛ��;LUs��&�8y��6,�ʿ� �,���i81	�_��_���-��$���@joq���'{��*[}A�F"��̚�i�N�������_�f�;��,R�1��vѶ����*E��~m��I�'�
��LS��i�� <��sqL��H�A�&W������Z䒐o�x��~�)��1V�~I�v�����|��t���l�pc6z	�Ґ:o�ӟ(K����E���F%%z���H}�u:P�L�����$ux�X�'�ͷ���uv/1CU����,���W�D1�<ע~�u�m� �Fc�/#By�Y�ۃ!����FƜq��S:��B�mv�s�9��G����^�6�4���\vO_��0/o��󮅕�����n�yz��)&�S����^��λ@�C��
RL�o���F'O6�MMà]���Y�4�oO̶��b�g��k�oH��]ir��#�m�Ԉǁ�d�xo���x��^��~�[9߈JE��V�_��4_n��T�f�6B��%��t����y?�2'��>�`S0PZ�;w+ȟE����/Ũ�W����H����,���:P2��$�/t����p"}��Y$�S���~�bu��2���'��f5���÷��]#��֟f�m����r�<���a4Qz���=EԖr� b��Q�2�%C�`C�.��>�8B�WȌm��M]�9�$�"�Z�.Vj��]�l�M���|��Q��'N��-���4��Wv��h��f�%lh��+L�_���}c���^��ir"���GV�)e#�O[��9|�"��ΐ�� o��x�^b/(��h|K�N��<�gjn�t������`� /W"c37��Zk��U*�N�q=���>��i(�ġ�Q�W�6���R�t;�'R̄vc��{=Tj�n�+hF��U�����.�J0�^̾8�@=)�P>X�7�G�H�rTJ��܎p�_n��L��A��2����ѱ4��~���X�cuF��<�*?�1�(���֩y�|ò�*6 �㙠�S�(n34?��U��It�m��/��Qv��X���Ζ[�W�|�T��h��Rq��vF��ydrʗ�&_��ޝ���7q(�4��)W��ّ�eiD5 9�&$�)����E�_c����|�	��whm�x�("r�mA�w  	�.΅��~���eΝ���,?1�S�$���U�Nҳ�Y���IW��:�j��u���_���M>��D�d�]9Y.f�A��q0��ކ�����/5 "�I��Cepб��VtW�q���ަ�|7�6lp	x(11�_^c;j)�diZp���JS��@g���G7��\X������
������*s���X�d\�E���*���i����S�}�<�q��} �)Ֆ����l��K ���~� �Uۈ͝w�1/�tD
��t���
Jv^��'fh�!���:�1o������H����y�!�H��c�Юym�ϵ���H1��<A���D���9�E�e"\��*j�����E+�;���=�G�ϕ�I�5��Mt��I�n��J�0F[vQ�o�7S�J�Y�ha����\�L��,��4<�z����v"J%5v0+�W&��vns�f~g6���}'����>��(Ӧ��/���JgEw�y�w6�E�}��*9X�$G�VǕ��8~o�Q�hIJ0��p;%�X����=��x֛� /�#��:� �����$����<�e����"�rU. ���JT|��;�tv��hu�-��1>A!�6���X^�԰_n������3�:S�����L:uC�^F!pa�� 2%j�ؤve�w��zLM���i`�E����x�x`��v�>͔�˗���$<g��n�i�3���a� ���:{4�)0b�a�AB�	�{gU��_��D�s�2��諺z�M���A��~�PQ�/*��y�{G��5q�q9�6�q���M��pt�4�iFo�2;���3D[��� �[6?�������H�E�)>l�jVdx
r���X
|p:��X�y�2�N}��dj>
��?��j<S�6�n}�'�Op���txc?�12�f˳9J��߲����C�b!-��c�9�\{�3�3{�]Bh���:KpD��Q�}Q[M6LI�W����>�d�1[�3`j�#�"q0�d���z���a\l��wr�%���9�3
z�4i؞Ǻ�2a֮v�}��#f$�<}51�,Ah(vC̖�I9 .�q;]�OX>�лԾ�YΕ�D�:�*$hK��|V�,���P��C�]��{�f?W,!���W*��w�$Gq�d}\�Ԭ�}b!�Y�o�����`c���@Mk^�p���.όf̟Ɛ$ٶ$Tl��y�zj�cL�.�����CRP��F��	�㡑2�25M�%Xcd �*�ɬ��4y=TQ�L�\͛�sθ�f�B� ��M����3�FH�F�E+kx�ֶYy���[}�aח�_��c$��vnHM��6�9�K`��4%yV��+�	��~�u�U��͐���2*��xxQ���|��H�����*t��!�ju�s�NH��v�rt�k��`����bU��U�D��h�'�-V�`c��p0R�<d�AC���f&j/��$A�(�u5.XY_�N=��X���}ˁhś*h�5K!��?���kb�X4��=s��3;Z���ǚ0��#���u� &	�oK����s�yigd�.[-��� ��K������ñrS#�T��.��k9���8T���ȳ#�5��l��ɓ�V�ӘC#� ��:�	���^�r��P��$�~/�	aeT�#�&��������y�񷘈����vv��q�S8��?T����R(|e�OZ*�	}#p|��1aQQ ޲�(S.�ӈ5�>��v������hX#��iJTԒ�L�9 ���\����{���O��.psd-�1��x�ލ��J^4���;`k4|Mu�L�(�B@`3B����!U� ̇�c�Lj\���m+�⍹{���K�	o�V�?͊��䈯�/�[��61��JƕBH	\�air(bޅ/�Ȋ��p;�w%�����z�7�E��:]�}�E�اPx����|d�Z�RnW��߱2"=��]��C�����h�MQ�0C#�\޹��	��Z]q�u�<SB�ר�ic���j�b�IV���{��M_.�Q���3�!��K�_��b���B1��h����}����ͷ�v�鲈<�~�S����9�P-3,'���k��r��
#�����壣��]�	:�T�DW�T>�-	6�@`(q�J'1y�����+��f�
�u�v�5��Akfշ�ŝ�)tM�3�g��gq�)��(2<�𳈂��2�����j2��5��K�����pґ��]<2�k8=������+���!I���pel\�س��u��K�;|��u��2�dz���Q1F����a���C6Zz�wq?ğ�ʪGr�9{�e��&{����݁��%���{Y�h(�J���_������W��x�P�>���˷d*��[׻�����G.���8����m5�e��)0��?�Ԟ�����]:�G�\E��`���X�ϟf:���g�..����k�t�
TAI1�1PX�٥B�x��@x�QA}LyI�l�M��C�G�H	=]m���{'@r�U��kΉSNu���d1돍^�uZ��&%�	�)�/�_�I�w��>b��<K�R�Q�7װH(�� Ѥ*=�/3����Y;�x��1Wŏ"fW��}=˘�F`��E�k��/+pA~�N��YGI�)�Q��00M�Y^m(v�w#`��������P��-\�?!n��Q����=���8�8ɄQ�3��qWy�b�K��S�C7��6\7�2A�V����"a�e�ɫt��:je�;l���:v���3c�D8�e�C%4�n��6,�K����)>�37�<��8�OY���f��ElK�lC�>�|J{!��g��N=�u#z�y��2��t����2�u��~r_2ˇ�7j��pX���F�A��g
@�ވ&��.�]Ԓ<�����b��[�#^�6�QtZa���|��,)`���*��
�W�r$�n�A�ʎS�X�,Y��Hn[��ǉd`������������|�Q�ۭ���/+ލy�V���?���/
�
�������ߗ1t 77�?�zo&i�mK��N��
h��\?
�m� �~#D�H�B�������v(�-�k�iQ�9M��vxS��4P֑�������6���p�\�[���������V�\��b��7a�aU/��6G�oiL�̶���ʋ.�4l1��e���U�w ��8��w�Eş˺�O��Bx���/�xYF����(x����M��p��!��|���z�3�	�[Ą�w���(g����?�M�y�����]�/�q�M�� a���Id/Ǌ<չ�U�H4���*�G�|ޔ5V�o7��2�Gv�?P4.��_�$\zl��
_�6��8k�5:Ʈ�Y-C���ds�~+4�*X��{�E���[&[բv<�62~���Jm��ؖj�C��ǅ����P~��>��?��U�p�6�9�c!�8δv�m��+���ZGgt{։a��^b:�HXpչ�.��1����h���z�O�uw ���d�]3�S�*%��{�m'W�d+tj���r뻣�"�ƸK��>;�>p��_Y��Ģ�X��6Rt'ʍ���Ь�Ƌ K� kG���0O�����S[v���_����
}���鷺�5Hp��/�3_����)Ͷ��� �=����	XR:��b��Gj�I�����&ݦ��?@v��۶U�i
����d���GK��C���|4.��|���Ea�����ìWV��7������1�ҽ�ҫ-����AYo9��(jUf���(##�@1pi�������v9�q
�I�M)�D��q1S������haPG�J�1l�=�}�T:�J�����Q�C]��^�.�A ��)��#9�Ν����wW��o�j�h��yؾae�����NpZ���|�`�x�̐̆0.��P�uM��%ߓ��_�n[{����;�z�~��"���$tj(���}s��D�ƀ�<��霷�&���Xp��l�����*����HW�@�w��W��dl�Ce��C�4x�ݢ�ͣ�|h�5�����*��:8j�͐�㻍��&�=<���ѿ���9��H�JTH3�F���4��	�6az%D��֣Lۃ��Æߣ16�jۧZ�<�n�yeP�:5��0M
&׏�H{w9K��� d�W2|.��Wi��>�22K@a����OvQnI�<����ݑ>�@mkj ���|B�'g�E��v�	(�����������-s��Z������IA�۲�ub>���Jű	��>p�C�tD�^{���8�8Z�/Õ�S����;.Īh��p�0�$����+���-�pB���B7ȖF�Ṣ���z�/��������Sy� 1�lƗ��t;*u{aƑ�����Tf�K���s��4S�c7��CW
�>�zV�����&􋩞a�^��_�V���h5��[·N�af��79$Df��+�SB�QgB?~�@��(�9G��'�4Z����y��k�pŵ=Б{]2�D�8aȦ�P(cMVƤ�/fݢ>.��Iܘ����Q0,��g#�����Y���\��M�PV'N=y��7~����8��b?����7��~:�`n!'%N�	�k�{!1���D�����_�[�R�Z�yL�����7jݚ}�}՞g�H�<���GO���*l����:D�l�:G�Y�3��`�;��v�8���қ��ء�O����7��;��Gu�~V?'�<��&Ǐ�)��>طd���0�XQ��)�	=W��3�=����t����}��H��/��l-����}�uzJU�}�N����cf��0 5��N=��3fX-2/��K��J!B�=����o�(�T��-�����3Y���lWE�
�&����c���j����-:�U���-|��^(�C8W.#�P���5g&4ҏOߦ #�H�L�V\nZح,��	��������w��f��դ�{�t��g&5��R&�^��ͥ�W34M����tQ���)�i>=w�3��3Pa�O������-�[h�c8��{I����u
 {����QŮv��׻p���Q����,�Ľ2y�C5�7a�Sib��SJ�Q~&!A�s�9K�����g���k�@�Ϫ�H��0�Z��@)��l�3�rQ��DGJ"Ge�r��yc����v���Aqõ��S<��o�����MOo8h�P$��Y�l������q��M��m@���k�Y�O���/~Q�Po�_/�A��{,�w���3����
 �G�h��/0."��|��#���kɯw�v�hFM�dOī����%�H����N�� p9��:�k�u̍^hr���dH��o�g�& Gs Ǳ�[�YWϿ�'����d�%c������.�òY ��#9���D9�H[��B}i�44��uTu�ovL'�cBj`PR�1'!m_
����D��H$ju���
�/��M��t�Ữ�s1�u,�ٓ-˾��,-��ď_y\�"+��P����};T���z��`*�fw���,y�W��W�JQ�=��4�$M(a�ӌ�,����D����'	�A��1x��1^K���B�̕M-ȁ�Ѝ��N��-�OÁ7��-���?���]��18�Ĩ��q>�ܽޚ[����+�*}7�&_E�xi盜�*E����i��e��>�%h?Z`��B���y��B
_��VJ!�8G�J�[ޞv��\��H_��C=P��mC��Icp^'T���3�b �x��&C��S�~�'y�Xc!�\��Q�@]M���.h��n昜���sE� �]�u���e�w��:,�?Rז�� ��/ʴo3'N�H���&�A���Mր��15\�F�eE`A-�ִZ�+��!oU�yd�9�H�7�:��n��b���p{o�Moe�"�t��Й9�c��mc�sϙ��R��@��ǳ� �ܥʦ5C`ߊ�8�=&B`����jH4�����/̓Eg��|(����-]�c\r�:��Ҳ����c'�V�3�s)�yb����6ѿ���{�������u\e��r
��%�R�Fw^��ˢ�2�"g�I"~���EP:�ֻ�=Hu�W�	�����P;ј�����&��uU�P$iQ�M��5lXs����?�>>e��	Bk�4L*N�2�-����̖��e�nѩN�!\�;����V�,��5p�/i�<!������ cH��N��b��o�X'˵��B�!H���'�'�-}��M���c5�9Q�nY��7����*��0PO�?����A��(��0g�S�sw(�}B���`!��D�f�ػ�4���/[%|۹��9 +��Q̲��'|�� l<������`�>:#�2/ɲy
����O��`+�$#o�UoQ�ށ&
�(�NӱHΫP��i��p,��P�?1=������p8�����qo��ڳ����
�D���{y�loO��y��ּP��=��u�������2���_^by/��H�xg�0��~s�]���%����cu����A+p��G"��w��ipE�xZ��xǔ���ٜ�X]��))���o��:u!��)�JB���{t�C�C7�u*�JpZ�ԃ90�_4���R�j�����r���V��
߁�V~]�o�Xj�?�Z[��W�z���g8���/4jGAb���M��Z7���d�tH�t�m��(�[*����ҹ�*��{>����&��gB�2͡����1�R�us�
���(2�ε�<�]i4~�s���R'I*�E��U3���+��X���Le�_����&�+$C�9�K�4V@�*7
�/�	��^�
ҧ���M���޴M`� V��!z�	c���c�66	���U��]�e�+e:Т2R��~B]�•�".˶A���Ҭ^�
*�YUh���"=���QlFP�{M��`jkt����p�'�I�	!�LMS�+N�<�=�}�b�)GՖ��Zd�y�F̂]�P'����W��@�M}�E�Z0��S�8ug椕�O�{��mjU�j��AP�1�����%�ݘ��,
�T]4�p�^K�O9n�	N�oL�e//��if\�{3�5�X6�q����ͥn�!v�m��1�Z� �й-�4�v+W���!�c�RK"PN�z(�hK� pӏ	���Ӆ�ԝ�����Ct�]?g�FA�a�Ȱ/wP7���E&^��a�`�M�1�w[����j���v�&����������Hjp����DjLs��{b��U�9�퓽s5Zؖ�(�&}��j����
��^J�3K3���D�1KP�ˊ�L�8�H�b0��PI؍��V#X 
eC�Q]|� _��2��k������)����J1���&�������nv:Mt�}� �P:2��X�ij#Ae�~N�,�[��B��k
ꂤ���#WG��ǃ�Si����!�]I4(�I���B�˯;�Z���P�.�La/wT�j|=�m�:�9\U�(u	,$�����ݚ8��+�tUaR����3h�~��
��JQ�yo���Kgb�i,=>H:ԙvK�DzԞ�ٗ	U!:M�Ʋ  2W��N� "0(�w�o���E��C�	)����)O�ؒ��wˋqgŒ�.I�qY9��6���蕞TUIq)1��c��3#foP���2�Y���K]ᴕ*2?۵Бc��a@���;� T5鞨���p�[to�����K�bY/��AxK�
 o	�mBB��I
�����oj
��g���cF��p��r�L��z& )�8�BL�x@65BN&�z���V�1��z��<@5DNQ���[Q� �Kh?UjM���+*3���_ξ��������N&<n=k�J�'9ScŃ�w�isC��%A}��ܝ�ʍ)���JfQG/��0��)y�V12��|�� �%HD*j/�8�y{�?Uˈ�(���B�w,�#lQ2�ׅ_@��o��t� �x�uݢ8$-�s%��k��<����?V%F�D�'����&�ia7� ��J�R𜁨TOvFn�o��Yu��Q���\�P{N	8���_F��h,�r��֝\M�VӘ�6$��\��[<�f�Y�=]�ڝ�[9Ʌ��u���JR��Ԓ�ݭ�S�EB�g�R!�T�c�m/3��+*����Y A{��v��9@aWQx.�K����&�s+�ӮG��y�#���;P��?��i\�kCY��66��Z��~��H@�F�3Ά�� ���*]��*�?F�Vg�5#7�rf|�/S��Bf��rHK��#���.v��m��O�AΥ�̽�Ei���ĿT�_£�dmOQ�Z��a��;��w�)j}tg�:A��ұ&�+�����E�f#r(��wq$�{��Ơ	�k�?����X;���'%����.On~���hR锤����P"<h��ta�j�}��]MWk��⯒�(���K�8��U+�R@.8��K{��;�\��T��؛��mZ��%W��?���\�#�pa!Y��><��D'�a���qeD�<�¦�G�A ����}�_$R5*�%�qm��=ݘL��A���g������O:{v�J�Uv-i���� ��{.���Z�n��1�K��Ui;�o�'۶�Z�w���'�]
�\�t7�9�R"���A	n�5����AonOz��<��;]뿊�
�B�?W@�}S�� ����+�C�JS�5��&G�eΗ�ڻ�n��-"��\I ���Z^�!�>�����CiL�	M�x�����,��}��ӂ�F�k�;���O 9\]�+6����\Z�c�j#�&��0=���ʘ��}D���?����H�V���SNZh�8#���M�p���%�sfկ���3�Ko�l#�w�W>��VW�f1��"��l��.�����d,����ck�H�!��wM�/tO<pF/�Ļ��$�D��ذmw��]jN��ڟ/]:��2C|�1��o]��<K�	25�ꉠ�pш d��C�:�mޓ�r�*�l�Y���}8�f��=��A���CZ��M�]�e扴|�bs�>��)lE;9��xfLS��=&���>��u�W A���a��s���!�S ���(�g�a��G���\~��n��=�k���c83�����u�r/a�S�mw�O��ە�1��h �ܝ�/�9X�ÈP�w/-$�T�=��f���b���n���z�x�F��%�����w]$I�y�~���vL�<�;.�Vzo/�"����ZLz�)��<[OΚl��ڤ��	?8��0W��h"2��)b4�u0^>�"|n�����Å6�`a�Sݐ�ȳ<��������$�Ֆ�@CA�N,�w���?m7�����է�y��'�0�wB�(��=;-L�,��zWc�pa�涕q���M{��������*=�����m�c��M�o�K'�:��s�ku�kЀ�̃�zwX�8 ��EgώV~[�`�'��.��m\��݅_BGf����Q�^x���t��[a�ѓb��&��Ͳ�o�"��t�uH�瀢 ����0��e�����q,�)�7�"���ţp�a���)]?K�h��~L�z8�Z�,If5��P�J��s4��X��O4��b�������[dmf����F����{G��*���x(�T�l�N[�g�3k��̘�h�4
�M���p�7ԁ�Ej�q"���`��#�{҈2
����N��*b��#���Q66�𱛪�f��v���m��<�%��8���+�O@�%E�I?=3� _(�1<_�gJ8�&�r�P�E�-{Xg�5�a$}~i�/��j~�a۽�K�X��	����[Rr d���~HL\��타�[9�E�5���"_*�Yk�8�t�E��2'c'��r����u�y��6��|�u�k�����2G�F�p�U�Oǣ	��>���G0{)���g���L����F����N!�H�<$D�0�ܑ0A$�U��v6�d�F�,�����g�v�$"������C3�[�~��M�we�1��;,�~�m�h�G�"�)��[9wh��
�@�|�d�P�����(]D��B�лM8� K`�=(@Iw���o��P�]'���M����2�^HT�
�`�D��&]R����Fqa|� �6K���?4ۆ�쯝�����PX�i�]����1[��unJ	�¾��������@=�s�TN�r�:�/h���t}��/�H�����I|��HF(%�\���	D�Ο��4��d���Kd���#�5݄�_'���ګpJk��"�@���֥��P�\�1�fi�I�\�
�T:�7�q�R�Ơ������3�
�� s��9�E
�UJH?
�/_ྟ-ߦ��|�r�ӂ$�����i�ޢJ���X�`�'�|���|��hG��e����y��br��;�&�ڋ[�p��Qqv�5 �)������"��{B}MP�z��}@��Ȱ.��{,����tb&�4x<H�k�z/���/��G�{��X*NBz|��(tC̽��2�����/Ng���j���g� �u	�9�tܮ�d�d����3�:ǌ���3?m��Z���T��5G���^�@�f"2�h�L=���]��˨˓a[ču�s�i��W7A��]R�Ry�#�P�y�>�͙_��*acO�'}�s���ӂ���Hw'l �d�d�<!N)y��"훀����/�����3�*�NVj��O����'h�)��:�S
�K��ɿ�@&�&�oE��b�V!r&�i�`Y�t4�Pz��:9���AڌޠI�,���tA���� 4Ү�f�Z˕ז[ϽLB��kG7����C9��Dj�0�fx�s��L�j|��I�A2=���R��)2i��4Z����B$��i;�
 �C�Jm/��f�d��%�zǀ��ك@=��Qq}VT*.�0��&5��+A��)k�r&�NL��?�n�n����i�?5�i.�yw�Ԣ'�'�v,�SbڊX�_�}���ޭ�Y�1 ⾁ِ�"c�*n;���p*���MЎd�h/+0�A��C�|�������j
��
�F�n^VK]2�eG�8��H4�)� )�S� *.f5�]<g 4�С\z�H��tS���� �-� C1�P)���\��w|ة�&�Z
�b��䱧r{�;��hY�xY[t����@��f� ^39�������'�����B��Ū.O1�7j�9lbv�kGm7��3B抔���b���*����ra~4�7(0u�f����y��Fވ�]S����gO�{��,���g:ZH@�3���l�L,��lܩ��v���.$=۷�n�s}(�խ@6�ݐB]����q�{���;�z�&��s����A;�,�,�n3������B���	�����1)�QUlb�x�Qq����9�n�	�����uZ��#����|�P��&+No�d����ctĒS�^�T�h�[�I�R��r${���,A��pŞU%R:bI�">˭��ޞ�[��aq�U������s\�Z�E��P �'�{����z�8��u5�.�q*��M�Y=f���SRե�Ħ׵����N/��D�@��=m͸1	Xt�ɭۊ�2͝q�r5�N��x|�b�D��L��eJ�5</PZ}"��*�5Q��re/�T	P�d纇�Qy3��4��X[>��.�>��`�������0H�9�4�PV�/Է��{�;�E6�(�]*	�w�TMZKR�{�N6oE�1RU/$G;Ì��F_7��^6��j-�7z噽��+1�r���#�Ka�e��L����׼�H�J���d�}+�v z�Ed���R]h��kP�	!x�O���$	���E�Ȩ(�+l9�hL0�G��Q��G�A�*gϮ����w��BᡵlK�/�~��*][��������84l[{����nSr���fԲR�ԉ�f(md����td�2��Q60�`�qs�ݏ�$�-w@]��1�f2y'�"01����-��R�M5��۠'z(�wIҩa3s�Kh˾�S��6���h��f�|�7�[��_�(e�,/�H ��°,�E.�w$�a�:`ݙ=d��`�F:�C,�f��Iu�2�����B��Ӯ�2��!�
P�@-��R�?�r���f�72k_/ݕkΥ�O�dG�;d<Q�=,�B]��%� Ͳ��-�=Z����$~�)R(�}��/����۬����4�A��h}ح��8ںjd���-w-M�\4�������z5_�����W
�#m��7�W�� 	U"ȅU�=�~[#<�؅b��x�d�lF����6�N�C���q&�\6�t��i����!E���cS��nq��I��z-u��f�dJ���s0m��-1���8N�V0km0���$�@ r�M��7�_L�[� T)�T��}&�j�w��{�3�^����l;��V���J�f���^D���
ޜ����*/m����!�X�y�2N�i�Y����xO4g*�69lO�I�Ȝ�LƬS�Y3�]�7� ����v�pM�X����\��T1���0�ʴ��Tt�����V�2C@�C�Db��icZW/�WX�vz��O��'�䳷ScOLA��ɲ�(��Y��<UA]�Jٶof�jދN��i�~ 7��{ݏ�Y)�XT�	�f�jW��H) Cdf�aD��҄�%���g����SL��p����3ҕ��m�$���a�����O�0.�~Z����2>�K�� Ӏ	P¹l��H��
#��G�W6|�-BV��������7��0$�"�Y*��9/���
�Zx	?��EҽSRʸ#?PsF��h��[cj��@Y���ڽ�ίnV[EF!�>�	��^�^9Y>\ܥ`$`�R�nZ�:`����MFQ.����Ĺ�:��!֔����)Xu����Fa�n�(�|\�<i�9����t1��d^�@�ɱDiU�KH�C�T�R�������M�8[y�kr�]����f�Ǌ�� ���>U~ t�e�d������#��zL�W6�k��u��|>��y��D���kZ�7�6�`�[��QSZ�-/�gSՋ��֥��:H+F,c;c�T���2yi�Z�v��Ai3Yy�x�ڳ>�#�G�<�E��%w��dp�X���H7����u����*VuLVP��x3����zV!��GB[�.^'v��z�^�v:��@�*���[؆b����2��Us���L^�+ibc�nHh5�d����u��h�<��5)f=ڸ���r���dK!��U�k.��^��u�k�G���~zhrU�m1�v|��ƽ��fp��y1U�Z��b-*�~hB�Ou�f2��x@�%�h�3̾�1A�:i�6�Vl8�����=�^�c)fl��ˆyn�USh�ە���w;UB���$�B�G����f�3�'�@���$��]��t�+�\���7���}�/�c��S���lPl����y~3���)���뉽uD�m��3�-�=�*���E�Mv�.M��ο�N��6Yi[�_���~����jT�x������oG�������أ���O��%m�^`���$!��a$ɑ�ǜ���my%g�is��m(>����g|�Y�������5�ʔ���\��R���K(�b�3��� W�_�0Q.Ŗ�t/9�؟��/�F`��gb\�DUqw*1�����1N����n&�"^��v�����YE�C|�I��=ٍ���&�Pk���*�	�S\�`ӕ�b���7�MPr�M���/�z?���I���V��2���� �����e�lV�C�v,�E`�"/X���g�?�zU,I��$��$U�<W�OY\��L&mP�}`Px�DOv�R�^���2I��'��L ,T�3I	�"��ԌE�8�/C�P�|ȇ�/ ��n�Խ�	F/�A�ig���ϋ�NlZ
Z��t.�=�f���l��&������?��.Ȉ.a,�Ug�5�҂���cWGu����:q�~v�!)y�<]0��XR�\�VHדT��:�em�\v�Ր���ٔfer��,F�w������7��uz�>J˳�4>�_�%;�X��V&;@��r�g��zE����eؓ�&��������`Y�.���/fg)I���#Rj�d��[6����,z�n��`���}n��hb��~�#J.塅D�ѿ��Ҿ)\��7bu*x)����-�j`�<�2�Y�Q��T�'ɒ(�]���1ͻ�]�:i)��Kʵ#9��w4HL۶��f�t0�v��M�0�]g(X����!
�.Z�kg�-��*+��i��C�U� p�,ۯ�H�*]sz<h��Cm�H��5{�Uʙ4�ۇ�"���V�P�l�S �����C�#c&�HJN.	��$�`y�fiu︀żc��>���|up���M��5q:�z=Dt��GkE�5�"�tj�_T�ݱ+��Lk+�5�$H��I�&�ﺂv�[��I��Q�_��6���5:b�~��+�w�M .��5ݴ�c�I�Dn�ν̿��O������P�S}"@�����&a�K���#����/<Lb�7��_;4�FoxE��rzu�?7����5/�D�Dq7��&�O7�����Dhemo�|Ǉk]Ⱦ�gfv�,����EV�ɷ����, ��aN�2S��:����
���R�3��M�1f����lʎ�wf��_��XJ����Hr�����h�P��$IRx�[ ��j=��7	�}Դ'��� O�a�M���
>֧Qb���X�+����2f!�u�#Ea��I�m���/n4;P���k�[	�lBn��p��˄�����\�E��(��k^�e��'�m7$��:P|�_tQ*te>�W1t���A��S�_�J��]Zƌ�&��6h�گ�7�0�b����(��ԓ���M��������̼ަݢ�,'��5����te��i
bť,.�]��$���p!��b��`C��Y2��doF]P�Th�]Wd�eq�����B�Z�/`���5�Q�8�Z-"�Ri	�w�yE�e��9��-���{T/;(X� �LgL^�w�3B�8yG��a=�s�]� ҈(�c��p��g5�H��\e��1�s���cuRqw��c0b[�\�^�Gx�UK,[�������z�)\�~��d�Gu`��	0ݍٿ�6 �TvM���`}�芉G�@S���}%�=��$��?��-!R*�����>�`l��8��]J�*�����CY�� 8fO8�P�[��کG�囀m�*+E�����p��IbRl�=f4�`d�Vu�>�=ӡw3���ƣ�5AYH*�Ne�n��������A=��d)��̨2��<���}�T��f$4ΔlF����r>�#���ã�.�m�k^����(8r�X���#�7���r9
�4�*�ظ�j4'!�.���EZ|�'��p��紛Ȧ3W���U�&�֭ �+�s�Ϧ�w�=���L�0!�(I$��]�&1fI���:sD,\�%���l�ibŐ xU9���3�ń2PPL����d��/�� ���2b��C�kU��TJ���T�D�I:0D���<�5�����s9\ ��/��Q?�cݥi7݌���<�h���n0��g�Go�U���z~�<0̯j�&��tU&���S���'e��BہJW{� o��L�e�6m>b�}��tJ�|����G^(U��[G&�`��RI�*<d�9��?�̟���ir���IIU�4ߢ�%A��5�n�;���ss�b|�N9��4�<���ʴ��߇�?<�� ������s��P�:�~p��u�Ƞs��Ń�HUI�9N�Q������@pP��F����m���w��ha�iEe�xo�����zy��E��&uV��Q��J�8�~S�����#Q�ͭ�ƫ~�D��ϟZ� +ŬJj��S[ⴐO^C]��R�����+ ��NL�O@v�����D|f�k<--L��y�{��i܅u�,AS��Z��$s
}�@л�O\7-��P���|ST�y�������$�e;-\��3Bd�\����K�Q�юO�g瓒�d�P��EY��(�uq�>��1Kc}��X%�Z�r���GgQ7u7� � �S�m���Ch�`���o�#��ƞuv�32���O����HNE�Fk- pT������Ӿ�0!.��dNV�X�N3_Uߪ3$%!&�<H��ɠ�{"��MA�|_C>��;?V��q�Up{)����%��Jq�%�hp���j�� (l�Ph��?M���H�!<c\v� ��R��2jS�g𨴔�A�L���{7z�\���j;-4��|��.{�^���_��'>�������Lt^5���!���@����[Y�)�w��z�a��E
ސ�z% (���˖O����Y�#�Nֳ�7�U�(�Q��mVOb#���F�S9���^~؃��Ԣȱ7�➄L)����h��w��~���7�Q��(��Ԇ���6Q��>�!��ϠA�{Մ�e���1����`�����<ƫfߐ=:�-�b>M��E�f��@�om�|,)���m�5L�&=+�k���=m�b���!X��zc�m٪w>&���l�PH����)��MA�A�m��ˆ4E �����q�4}���-�*Wd�땉��0��&.�%}�D};��������20�Zu���
��J���xe��B��F֜�up+|�/���Omab�a B�A�k��w/"#*��_�+.��ȉ�;�M�E�tA�#�w�z:�0O�0Tjvh��5j�A��XG`]�|$GD��Eu�����#�q�!w��P蒎����1=HS��&+\~��X ��d������a�/��̰d�u{����oa�.1��7�����Sx�M/\����ȸWb� U��=��u�@��͑�a|����`L ���uyY����:|C�g�BE#w5�çP�y���}��.X�D�Z���m��Xn
��1UAB=�지c,�5�f+�>YV����~U��o��&JV�����h�� B5�_��k�sr��{�*���~�v�b ���R�i�ԁ�^�|f�:��xո��4u�);�st.���F��&�&�0�@@:�0J�H���jE&�3�" ������78�u��U���A�����k����P�b�����'�����bQ�b܏U:m0.����@Qц�yw������F�)�dN��}����^�D��$�W������dI������B ��w�_��V�f֌["�H=���L�NfR�<[�N8��w���~�Wܬh�rFPק>��1_ ��)�5������N���P�Y���*[�ay)8��i#i�Qx�蒌��@H�!�x�q�1�D]+��ťAߟE��H')�1I磠8��M3���G��t2FQ���	������ŗm}�8Ռ��GN��G�Q�8��f_���A�4$>9���0<THM&5�ϔ�oi��K{q/��2W������9؊*�d%��
�̹N-��8�N��O��D�^u�Z�:�"Ҁ�Ƃ;/�©Sv��e�<��lȫ̖�#��Hۧ��;��޽�r�_25��{D^g��κ��f�z�xÀoy�����LޗaP�_8w3����ZO������O�yw8{��xw�Q�1�0L����@m>�[U�0�+O��3�&���
���+�U*��
�n�!TS:�XT������`��3�����[�I���l���=Q���P���s3��Q:Bȇ��Q�ܯ"��j�G��߰
Ǵnq�|�{����|��s�Ո�*�B	�5��KIBm4�V<$֧ź�0�a��Ne8��-P��ِKB�+���dGN&��#�j�X�@�o1K0���`�7�
;:C)���Ȍ����b��ώ��T�^8s<YF���iK�h^ۄלq���q����-z�o}��=H�+�&g	�����kw��j�[!GFw�骳;+y�I�8��kI�.��-�M�2��n��iw���!�~T�;�tJTjC|)E��g��΀����I��7P��a�d۾�P�)��ߦ�J�g�Z�Ѧ�bu��Q�XA�@q��<#^�A��|���ȷ9ۊ_,qE��`�.�H����5"3���ބ�M\ s��P�L�����"�V��Ք;2�2�AF����x��e]?Yo��^-�F�
���.��٧X���u��9��\�j��"a`��u%�`訤��{Ii�г�Շ��!9Pu�8E�4D2�pۑ�tRj�Dfi��;`�q����$��/�E���͢Ѐ��
M��x�B�v�˅��� �v�b���Kf��s��Xa����9�D�aĤ�#��O=&;�9�m�~c���x,�)B(h��d��oy>r�̶w����R��}G�f� MO#mE#b�iˤ�R�e��P �n]*��Ua�]'�� 6�O�;18�/���<��u
�j+���&��_ �t��EB�T�?����m��c���X�܋�̨Oq�O������t��#2���t}�Fj�^����u��շM��m�����aQ*�w<��0��~ ��1?r\�w���*��G:����9|��p�IT���-�<Q��xղ3�gqb��������p���N�1�sW�q�� 0�<F�#L��E2�� ���u�'��`��J�tN��{7J
�Ѷ��WD���rmg=��m�o2]��jiu�3X��O�i����z�6u4i�C9�ZZ�_��v���?�&��ru��r�d�?Rt|V���Y���>�
{�O^�_�_�3!�í0�F1i>��
~O���wS	�m ~LXA��9�#��'�c�ˋ͆V���d��`��գ�&FB���5����a܂�lJK?���"���Ib�?�/IR��gQꁋDW,|��d-]C4-�D�,��vl��Y���x �&��1 6N+�C`�)���vS~xIU�鬉:����ӣ�"_^���zq�zbg>,�� /C�b�'_[�e;wD��`���a�z"�sɾqPU�d����؈�u:���0fOu=>��HѳI�D(���7�t�o�ǆ����H�Ҫ�9v��l���>�-�X����5��8<J����P���M���K�a�I�Vq4�:6�s�h>�o�����a��I��&�r�C��c3Z9�@w��rٔeH#���Y`g�K;3��3�\�֮!����Őt�	^d�%��e�|�J��E?��J�k�R���s��!�-H3/�Q��f9��af7;1A��^��$#|�z�i�D��wXE�(X��ۻ[տ�zx!갋G�aQ?h�e����97�������hQ<g���A���G2�7z*�m_c͎��3R��j�N�ݚ��<SXq'F*�x$�a�=t� t~HA�'_�^s�~G϶T>�G�{`J�v�ǡ�W����#l�ۑ�ROh�O.AH�=�������yC�|e�_[�<˲���>�-Y���p�CoVyN%t����ge��HZl�F��>�H��J��������ͪq��/X�wIGN�D��~����O�Sh���֒��&"o�9c��)齁���*��	Q��{�,%�ay��X6 �܀���Bb%��a�Fэ��I���XH������l�;n�����]X�#Ϫ�,�h�ϡ���E�j�ܑ��6����Z��s���M(<�3�W~;9�e����2GH<�MT� K� 3B���^}��GE��R�(Û��'h)�)S��#�d9<�ۭ0S�>d��*�h�H?t|e͎���*Q�t�[54�Rd�q�@��|V�;Th�8i�g��)EYշlC��85��Nc��am=<���';fKC� 0��?6_�����?�;[RY�e�s	3�K�#1c�A8T+� �����ڲ�[���I��	�qX�5�vəEк�\=&sG���	��_�年\W$��W�)LF��;�02bedo�� _@�B��
��i��gu���27�b��g�x�wX���v�~K\��ߩ �w��	��ClQ&.��-\�f��4����h�����r��Ͱ�N�����k��GH.�~7[P�{��y��cgg
�hsP����-��z��eM�Ff�`1�O��j�2�(�e������C��w�PJ�?y~����8�xb�G��"|���LcK�xQrh�'�Sa�"�Eɓw? q�%��A�`Y�/��;!��JM��A��uvq�	�G���O��Sj�Z\��P�ރܤ8�>Cy��Ӱ����P�+���{vB�K�iec�a�A��+�P�8a�y2�Z��&����C;�[k�����>���Zq��y��3`C]_>�-'�:N}�=T�C͎��/dT6������z�&���<���A2(��q�"����1��\�B��Q��&~f��	��<����na�<	�����]c��;�2)]/� �8k��sƘ_RoV�D/� ����$����N�n*!X�פ4�ΖU�Q��;�� ��n�����yF,	�����`�^�S��@�jЫŷ2�]���#23�^��*�`�n���mW�<b�bkk��;5�Y���6���-ޯ���j���@z�Ss��o?HV�:@�o��x@W;�֡?���?��&�7Pٖz��v�� !8"rO2��mf=��"�n�\�<�Pj���d�Ǥ�x�P�=�nh�H2/����dY��^&Eb�u�	DN�!soC*�uU�_ I��2ظ�D�OѰ�Dx����v��#�$�/��p�L>xw�t�ix3�t�ڳuk`|�; ��a��pBd_�)K�pQ��O:���uQn�n�J6;�,������i�މ�U��������m�S�E���uQ��DLBT/��\�<\�
���-C�hZ5�$?�	�ϾC�5�����$\��u@�"�����T"�B���ϑڎ%�m����Q�?�z���x~��s�.��$9���j,��$�H\�J��Ki2����������|f�&�