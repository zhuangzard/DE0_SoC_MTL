��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d�v<��m���X#�m�o*�����z5�22�8�G4�x�{[��IW��(X(_<A�&��աW��'�mҳ�۫xv�<��
�5O���q��z*�\�"�ł}ʙF[BT�8����f���Qq��A�?kQ����#���pN^�}�2P��3�;��UD��UVҪ��Ǟ�H� �a�C��|�� �P�'Ђ�����|o�]1��%���L��a�B�JN���9�k���yEoȈ Xͬ���j���*��y"F��Z�G�>�FR�+�j�*��u"�pސz�x�Z&<�x����.s���r����.�,��0F�a
��$<&�s*K׵�����G%����c�܇,Ŗ|*�~�;ɹ�z����$���w%���{��`'���>���h�b3 X/ұ�Z6�@�úe#ә�~R5���ïSQ�C�vt���= ��9�º>��F�
�7k���4	���]>������ L�>��Kh�{ꤊJ�K�\%Մ��E�R��>�)�w�c��;w����[�啊�9e��F�|�$䵜,D��-e��6p.7���g����a@�UYl��p�������q��eS"����+UdM'�53= }��q�پ�I Gq")�`j_i�s%�%�7r-�G/��&D'���ԫ��a(�bX1Q1�����7p�6��x9��B6@2��i}$��-�n���m���3�/��DG�M���c��~dۮݕ�rja��ѭ�<�{�3f�n||���q`�3��u��^��%4�:=?�S���π/t?�B�j�*�=F��
_|�J}$q�)b�W�(.�1P��Q���T­+�|Ω~�0,�7)��L+ځ���T8�8�$:�����[J�0�<�����K#�E�L��J��e��� ���g��G�5��X���:5p7�+@X��6�N��E˸΢�G�٥`{e�`z���%D��8=���.�.(�LTlG��1���IF�G�A����XzY�H}w0���wh����V�!b<�����k�Rwn�H�:,�=�����ՠե5M������4o�#i���=��҉�
���57�".�-3��%�$��Nx�i����Q���������``i���w��L�&���������q��D:�>�<*�TJ+�V�,����	��մ�0�Zm��U5*��W�@餎\�s�Nd�z��/�P�_j��)�*Ja3���_ߖ�����ī�r��Ų��P�q��R���Ӣ��	Ng���+^��^f�#�l�S`�z�¬�1�{�7��$X�������m����tx3�5J#J=�7�a[�C�H5C~S� g��_� ݔ��b��8���}�6�g2y����i#�)���#�V.��\9��{��D�/v��[?����B�,��+@��9N�5=��.V�0����mgH��'m������Gj�؟��5DeS���R�g�Z�OC� 9�}ބ��*r��2��O.e<r59m�= �s�觇��ǃ*�\�P�7c��9�1_�ކ�d�yE��?c��\ƞ�c:^�_H�S�+ɽ���s�W�y��TM�Wb�1�7d��o��.��a"��}Vp<���Ⱥ�Vb�h����P��y�.�	S�ٗ뛟��9�"|Ư��@�9����ei�g�(,�Wz �>�*$�V��#�ڗ��g����5�!�E��K�ֈۋ�Oo���A�$[��Z���|et1\$��R�j�1��5}B����$�m-I�6��]����mљ?氓g���o�Eot-����y-���jӂİ�Y�����ƿ���F6%�w"98��UHU{��v$���ol1[4��I��N�e��݇�������k�&�[J��8�wDH��8-�OeW(�lMȢ��Z�҉��%��}ɞ�K4�%�E�S��^'���?S��)z.[��E���{ij�:	ځ��.෪"̈i�3�a�tpY�PVlP�K	��EL,=PV��3����M�d�<*0�T�G�ߗ`���i=�F�^A�g�M�b��d���s}t���>M���w��W�y�f*n#"�sMTG��;QA�S*��kQ6��G��\ �aс�,�f���b�����+7>���.��?MfXn˗�Wh����T�Tm��������pW8�'$�pp��n?���>D��������_�ea��~��CbJ��� ��0�uM�u�սn:���2�V
Rd�;�@�]���n�����]z糞���F~���趀�ǪZ
�lڲ]�n�WE
�@?�ǧ�0��![�0 �} �^X+g��>��l�qL��>M���5;1�O��BQRWfG�Q�|��I�O:ǩ���w!n�焜��&l5q��?!H��V�:���%��5	��z|���k��jB�$�Q�e'� !�i�Hq��ީu� � K
Ȅ���L�&�ckW�k&"�Bx�5g]��'|;{r�)�n=�|IK�V��v�'�������� ��<��^��2C�_���r�Dg!�舖J��^Ѥ��\:o(�\�t+�����Z[��6�S��_��8[��"��x}�{���:6$�YB�L��+���+�&35��R�rqvB�I�}J���� ����7x�\n3=�IKǰ�`じ-?��x�\�����P;����\h�_����vM]�:O9*�UIwX��ïKqA�c�.�:{�=�}c�'�S^���X޿,����=�U6EC>m }����q݂6Z��`�p/�\��\XA��[��5̖}̊a����hA��s�k����Cb3�)�,�\���g�� �ķ�`�I˭��hei� �b��&������t�~t|Gq�_�8GF���A��q����E�E�/�Nq/^���F,�JhYN�+c�d�f���x�u�_k��q���S��qX�dI
��H�c���y������	&����4�����-"���=l2
Yb�U����5*���6N@"�@)�,
���~?;�wo`��?�hf*�'�Av�:���2�X�= T8g[p$+���sCL8�{ 򃥷��2!W�!���@%x�]69�c�2ܘG��Y�>����3��WFI�����p	� Ƀ������I�o���!���|�~1���Bes�e.���"K�>t��:�ɱ��&��+t�4B�b4hH���وQ��ZaH���+WH��4�T
� �$��<����Ͻ�Zc|����=��	>����-���L��0JS��w�'z�%]�O��/��A�F�[bbr�5��^Q.TU���ek')��j�
9l��
G����#Z���ʔ]���'<��o���AT��0���J:�^~���.�*�ES�ȓ�9q�[oB6�;�F�[�l����/C6��g�d�;\�81��x�Ե���L)[,z �+�i(tan���q�o#�ׂ�-��9��ZOD-�_��zڤ�w�.{�q�n(X,/՘V��M#�l\��@WU^�Vi��Nl�Á�r������@�+_�R�n�NdD�Ж.(���3g9�j^^!-��|s����~�s��[!!�Q]�-�'��?�.��|��{7���/�r?��� K$?%PA�5����'�ݓ�E�	�e��|���3��k2h8mJTN�k�/�W^ %��[D�ŞH��r�3:����adc5� Z�Ш�ö[H������ܓ�}���^J�S�c�N��Ӧgb��_���~�޼����l�cx���u��S@W��:J�d@�y	�����$�v��&I�&�+?~I?_}���5�#�5>%�6��N�[�8m*�����H�4��~���߼D�`�'�n��ZPh��b+d�b��J|����Ki	< ��Xq���}�ۈ����Q7�`��%�\�-T�Cɤ��QOɵ�j�A�ɸTHx�4�b?n@e�
%�^��IZ��Y�|�S�p���8��i'����g=R.h�ho��M�߆8M�gNfI�;��!�/�]^l�M w/�o{�̱9��h�C��1^�|q�I�'���R� �ݝ��zoy�9�����c� ��Q��a��,�t��lN	���qZ=�%��I<������aIzĜ��Ɖ7��\��J�3W;�������1�))�j�K.7��w�'Tܾ��	'��%��V#��uI�� NH��F��Ǌ�n��:��[fDB�>���+b�Q Yt�,2�WZ_�������ư�����^������F�3t�C�����Ff�����	o�Y���g~kB�>��F�3�~�󩘒�{iP�iw����5���L��^�Js.y�&y!mu��foR���B4Na'�6x����xpv����X�p>�lR$������;�uT����@d',ڻ��;���.�����F��H�7������$���:$ZZn2�K��E��W�|���/(�GL kO��В�9�_�'�=׊���閁½�H�S�|?|�L8J@�G�3�y_E�2{"�C򥏎UsK�����F۟�D�|��Z����E�����)Q��\0}�4�;��$)��Tㅿa�M��������hQ�	����o�o�r����%&�a�(]�b�#nB�C�Ѹ	�>�R��`/U�a�gx˒�/�����|�㋒�Ϡ�X��S�Zpw��m����p�]�yH�+��MD�LB���1�5�|*u�Lzn�X�<7��wg*���?����kf���3��L+�)�}v?���������{r���^�NE��b-�͞^�M���O|���G6uB �uߋ�%މu�C��)��zT���ɖ��tU�-E&�5�o͞eM��&��eoG��Rw�~� �Uob��Ċ�@���V�Ppi��q�a�vg"݂�1'�k�wC���dFED
��Y��'~e���4��J,Mp�A��/�m_��&<�(]-�Œ�@h廿
?�Uh�>�gm����7j-�ս�*²�?��m����;Qha��U5 :��:�&����Nz�b&d���[�$;��X�����(e�$citX8sB-4;D�#:�K''�^��i�[��Q=������n�D��cb���a��?�ۏ�ű���l%\Fj�~�rJX����u��E�@���P�Ȱ}��~�3�e	��^4,z�u��^��k��������1�����^d�<�T&��^��y)b���NOޣ�������J�/�.�'�g���}��@E��{��S�n5��-����Q�뽒�3�f�C���י�4�L���l=����Cu`Q��94H<���(:�?V��o�)_&l�;��6JuA Ol޺ �%��S��Y'x;	c���=�����k�̺�+1(��;U�";R7Ȯ-p���F����2���k�2H?�V�G6V�gC�WK$>J���#���H۹?��@Ӝ�+��G�vd�K�a�kE]��Xܢĵ�M@�.�
��®c�����G��Z��,��,>3S��E��>/tw��-��ɧY��_R��ss�o5w�Ta /������4�Y٘�-�2ɡsh�����h� �1h.,�|#�G��ٛ.;>tw�gǃLE�[���#Rù�8�����u�д����	�XT����i�?��$po��^���<���%����pί.,�\5%�[�C��.���.-�oMr��l:/�~u����8�o�	ǎe?J�:1����0}G4l�@���yN���w.�;�Un*��n�����m���FX�⪪Zf5|`a_��5��M���b���8ij]HB�i�hL���-�B%TY���O����3��ԉG"� N�0_㠟�o��G��yi$.��פL�,p�K^�nH���K��y���W����>{rrt8capʿjk��x���xV�ʺn ��\uB��Q�K�R�����4��@Bχ���x�[��V��w�~��^=t��]t<��E+n`�N!��K�J*�Q~�NT�A���(�#�O荙g�<XW�[J����.!�B9|�,cvM��֚f��Xo��A�t���n�wU����~�J��l0��Qs��宖>��2��������n����V0�F� ;5�k�U�.�'2:�������kG[|UvQ@K՛�`���3&#�e�J��	2�"��Z��J�������w*�p���j��uP#Z��� ��W���*n��,�xIo�80�̜��Y{V��%٥S��Ri����ݝ\	܋}�sC^����d1E��s!�{.#60�u��p�Z�j�ss��Yh^/�:\�s�M�:���¶��NE ����7��!�^��\=N���O1�~���s.��{�3;^��d���8Q��:#���ΗvP�V%�=�ٷ�*��<3���#��!��J#��;�ٙ��I�Wf�$�6m��/�53:n�3~�IS2X��$A��e1M6.5]y������+���	���(ib:�x��ʵZ��#��u�zF��AV�j�i�6gM$i��-���0�r`�g����y;޸C���V^�#�7�Ѯ������T pg�w[5VuHq�9�����Ǟ�NB��!K������
��R5`��~$S.���Ë�+��	'��F`�5ԋ��2\��zs���8a,��u�J�(�y��Z���-X�����ط���ɮ���(��H0ؗ�獢ьtf�V��Ӭy�ů�(���X6 jw�Em|g?�@Y��hA�n�!��A,=�(G��jm:L��3��z� \HM3��U^'͏١]ڽOd�5#A��3U����kj�����"���"A�e�w!#-��e��)�ܳ�<O�C�vU�Q�u��pJ�yUx����4�j�ɴ�c�޽��%��x�E�D7���8���h+/�%���g�u�s��=/5�� ������*�|�4h�
�k��\z�M�1�@��"�y���f��!���Z\vNP�d��c�{��C�E��:%��4�x,l5�Cc��[4kI��U0o����� �Ͻ~B�L+(��IǮ4��K���!����д�0��>�.�L�V�6����N^b�	O���qp�9`��sy����l*�����f��R!�� �	L%�t1���G�� �u	��9(��!��G�{ 8���4Py"����*Y�����t���QaEJ7"��=Z��SF1�aї�훚��׿�Y��.�aݷ���܊a�h>l=3�P;A���%��~z�?���޻1�_}X������H�����+j�i��qg�vy�?9�s�GB���yJ�Y�̇�͐�{ n�ȃ���=��&~j4���;�-�G�����9Ӛ����mή	�����fR		�b6���n���9�����uB�̲�mlO'��R��~�g����I� �ۼA�+)]��U�=����]׃?�9IT��N�Q�3�E���9Pӭ2i�]��YG��&���Lr�!����.���E�/�����%�,9J����_u1f}»b�m�C�)�S3xbo�cGˬ�fR)/m?�6��(Y4[i ���#r!���,���?ᡄ�����$.�����yY4���H������;T�xS������n{ߓ����5�F��[����~��ʂk�аZ��רX2��G�*ƭH������.�F��lnO��yJ�\q^B)��@�¢�2n�k�V���)f��e�od�Q�]��ډ��wGz�h�f�l���L033q��9��S(��ϊTT-z���^��F�������󱛠M�)EB�鎠�ߙ;(�� i�9F|_;��I6n�E.��f��v�ڱD�Mg.�§5��oK:]DofAEqe���&ӫ*�g�Ѷ�p��������ܼ�a��Ϋ�l�v�Y3���B�����(�\�ڣd"�"?4G�>���d�"z�F�I6v��(�E=�Y�b�_6_ ��������g�	Aj8 dO����7K ���N�~�������9�GT0H��q�4,��,"���_	F�\���dR5>��﬑ha�Y�5����x"�����ux���\-��!)T�稄����%G�k*}fN����=�v�����QR��߰zD��9 Q��dj���;m{dp2��о#�1�Ѡ������H�	�|65���w���ROka1!��������	f^��,�@4N�V�6�K����n�!9�\B�6@#�n����6��SA��`�n�[(,�otP~-�/��.�����Wz�3�o�������qk_�Yn_�����b:GA��Ď�٭��B��l?&��1���u(�!O):y:���ٌ)�܌쥓k��mG˯<����lӐ��֥d�p��Qy��������;�������|�r�LF�p�v��6Ѩ3���O+��ټ����rW��x�AB%ZT���`nxoڶgU(��n3���࠶Y�h�@�PH�8�5D���J�U��Y���h��`c�  ��iHZ�98B6��������>ӍcS6}��ha��v�&1B�_��4�K��ż{��mn��]����4��o�#k�߳/7�q��H BdA.3񤷔���Ob⋏�R�a��GS����2V�3�8<��x�C��A*� W\`חvɁH��B�`n�����"��
��g������:(6O����>ɗ�S����!z8#1k�×D�S�����)�R5�A�U����o��(K�Q4�)I�Cg�	KX�����wM��b�+��W��A
98�V¯Lܞ�I�M�Up1jk�'�5!�	�/�-$d�����V0������;��0q[4!���F�
1���/d�b�����6�{flS�B�2�H}�M(��D6���}a^�q�<�=��V�"�Ə�ܙ��L;�*{���L�% |pg�F�����ofsi�N;��±���.	�.sE�~��:^�ۏ��I���g��<"�A@a�m�sq���=�t�����9��c��ak�g����2yF�r��0�ӵ���o�ʲ�O���c��1��-�)�bc����z{Ӛ@�^�d4،���[�&�1U.����+�3K{	$��{gˆdD.x����WZ���%
t����5-��ng���8�	_��G4EC�޴�|��>�m��C�s����%2Ж���3d��e�B���T^�iӇ!��W�Y����m[&Ʒ>Bg{��{����1�ہ��[uI���]i�ϐ��4ɻb6�`i�֟S��O�иd��"�M�\#g(4 �s�`.'�����&Z��~/SH�ٕ�X�s�T��Y����,��9S��L{�9|�������A>��A.��	8�����![��Ja��U�$���c�ؿ��%�h��$�����I��hó�U��8�H񠕀�ɦN������-���,�m���>���r��B���ͻ���&�oG{�B�-,mB9Z����'���z�9��Z�?MR�y�V�%��<N~v��~0 dؼq�0���<�1���f{l�Vf��P�AL�>�	�ϯ{Y�Ta����s�7ŀ�j��AC
u�v"������SGǊ]~c�a]�>��`1C�B:�H!C ��v��˒�u�PQ�]�ݯo3��Y�����t�����R���x��F��}񚂬(@�?l�����y����P�V%��&���XD�x��uVr���vr�*v�3D���� �H����DF�^M�-��K@Ghi�1��d-��Q������k����ݦ��f'�|3�S�=�m��.#XW�V@�w������@Р�t�g�R�?cꠇ�?ܵ�ꝷ{TBnP�\C���TRfj2m�0˧e��D��ʒ���%VM�V/ Y�鼄����N������Z �4�q�WSj��~,T�~��m�h"d�6@�����T�W�_�l�@aЀQ�%����=pԭ�}x���g�j�@��?�\ֳ�);Y�Sa�}e2ݲ�K���b��L� fs�Li�;�Q���Su%I	�h�ͅ9��Ỷ�	�0wl����R�Ԃ^���s5W;Q5ޙ�| to��r�o�ڞ��Ø��'$>������0:�)���QV��srw6Z�%���K���zV���6ݾ%ZL�A���b�ڍ�4�c����墇�����g
�;aL�+�/�e�0�h�x�g�O���@	֘�\�-�K�<OiI�i�¯�媺�(�H~#]�&�U\�u.L���g�}�\�nWh5�@-U[l��$�g�n�����T�|�*�����F��d�l���#t��n�%�8\��"}��G
��q���
�5�'�>�*��8��et�����|��|d	��>�^Q#'?R�s����ܘ�`��yb4sZ���,96-��5��<�QEP�Kz�� �#�Ȇ!]�
r�Ii(>��b+0[,VX=��|Ǘ�Á�]~����񺩊�a�����g���p���:��OR�q�4J�J,?l&��xӐ�|�3x�LT�~,���Ydku`�]�^�w?o�h�����Qإ+T��Q&���pD�H�>L�,ǸXZ�&1���������9M���+H��g�����&�sd|�%�˸��z�y�;�w@�kۛG/�Қ�ϯ��UH� O�~��\^�ࢳ���ni��is2�s���Fm�ٝ�TBƘ��p��bXi�խ�i27ݜ�5Dly��<�306;n�t���<�T��JX�h�GG�W0�k��f�ћ��Y돉�"�3q.��JLf��!�2a���͹}>w��Oi`���&�&�Y²���B3�U|�a�w��ɱ���S���%7�D���4�H�1�u�����aj?͝�]�_��e�aW~tdy�|���}4�7���|��@�	�z�r�rp�Uȴz�/1��X�电����@������Ɉ�^�Vw7��c������j|R�%�����S�md�DM'��[/�eùp�P��c��M�^/�K���12�\�L�!i�'������C��4\�����4�m!n�*�yfi�m^��Z�^j�z�����vqzsm"��DP�+h!�Z>?��	�|v�C�Gi�D�,V���n�|Gt��pK��,#��W"�O��'�u�t�{���kҼ�`[I5�)J?ЮyqC̎�(�,��@&���.�b$�TQ��S��F�Z_x�P���B�X@�Cl�c��&h�s�	n��)���ґ��e��}T��zs��
��̹�3������;<���fq0��XMb��C�b�����Nq�y�Gjb���S��?�G��)�7\�H�;�/�k���n)����U��P����d$
�"(�<i��z�U.��=f	`'і���{֪zONf6+D��X���N�5���k⧼`��f��ߢ�,��� �%!�U��t��oBݙyhL@��G�8F����)q �Z��8��XM����K�ppeOq�B/Qz7Y�h�Ŷ.gCП��Y�?��aK��|�p����3�W�^e���8�aU_��;wj���������	m���\~|5k1���U�桋�G��O��N�=���?����K`dea�f�U��u�=�7Q�ho��yç�!=�c?��tIV�KBӺ��cS
� T����\���{��ƥS7,R5�)�ټ��*�⼚�B"�2��1c�
���*�L Ձ���J�8~�7���r��8#��z��w:gz9ީ x'YEPD�iM�y�*�IA�/@�v��br���js�hM�ʵ��Q�P��di��ƙ�Ro`\J܍5��
��=o��oͫ���pHi�G�o��M9��ͧ��_��Y�wV͚�.��&J�ӿ^x?��_ږxhm��hBס��-�0u��?e1+��M��X'�r���wQ g?6����w�~<y����m��:�6��=��b�q �3�g���W�`,k=�-)���y�~�i����!�p� �X��FB/�u��}Wv�j���mw���g�<��Ӱ!;�.��O�>���i�NF�t����_d����fGU���?�3�Z'"��k�,��*���S�x�,�Z��^翰��woHox����- �l��kҚ	�	L�|0
�s�*��8ù�Y��*4��+m�B8L�P�p��D��?-"Â���˃�(�q& �A�"w��	 i5	�ll�LUx`n�8�����!���hpL����@k?NSy=�<+�ʰ-�a+
��]�j�A��F��%?����n�,��I�e����#t/�Ʃt��cb����J?��ęW$������*��'�r �m�S��$���R�\���-��C��J��&��W�t�fY�����s����P�!3 d@�5cSځ�\x}4��"ß��W'VɎ�j�"&2/�?��~�<3�n��r?���%�;�%_��Gk�>,�u��>����=ȝ	P��
�Z�����&��徒����������4Q�_��-�IS}�<�w����ے���.�z�Q!�ȳ� ��s���	�ܬ�)�h��v�'h��z�cos�k��ϊH�Dć9u�y�J3�J����^6�۽�pM����*��Ђ\p�I��x�_8��oL c�IF�Yw%���JCj����*�	��lY|�P��#0_%�ʃ[��989g)��C0{`0׹i�c��U�A��z�3��۪/B�"P=%���P�8K�?
�'/��&g�{�uP� M�U�7�}c{2B�	xK<���a�(D��>���c)�O�i���<D�n�[��;y�`4�Jl�}�7����/ߏ��Uƭ�1vi���k\0/*}g�
�L�C��a��Ҫ��,�D�:#�K�=�î���H�[J�����N�Ǹ;~���x����y�H%?,�(:Qf�h⢀jx/���5��Nk?С�	�Q���O���@�c'2�}��/"@
%�RI�$�fϷ'��O�� 8��Gx�خ(�4�l�8��/���6���GF�sWv�,��i����F���K*�$q?���1�o
R��m����x������$�����[����@�ɫg��AA@���, 16]�2Pk�Gqۄ�r��n/��n&t�$�f�"�� � h��-�5����oCC䍭;�}�Ь����sT}��Y�)�ϐ�+<�Bd�J�!��Tb�qШ���S��i+L:.�yEP<�1�1H\�#��͸�s%��.��xw,����Z�(��Y�͡���_G@b~䕣bV�WΔ�x��0z]�%@ۺ�j�?,������-�v�n&	��j�
|��W�&�|>b����^ː��]NS�R6e|���{���']�����վ�եV��J�bi�3���6p�Dԛ\�h��/�3�8���g��y�����)�wV�(r�z��F�!S
��C�g=tQ��hl�2��X�`d�N�r�OE��{f9�%�MR)}��Je���v���[�֑��J���k��&3��]��R�P�Q6<H3$(���x����?�q�G;��%��6�u,�p������<�Ŗż�v��,���Řz��e���pK��5�f��H�	���cV��:�3���d�Wy3 ��������aHF����>,0���Ѐ͜�Ceзb��xs�x�O3V�c*4�_�{76�����=�qJML���a<��o#BA�t\����a�J��a,��j�s.�r�?*���4p��G5:�w"���F�������5r)��M�C�����{L�R[�|s!�w{<���\��M�7LԢE����(�[����S���!��]G>�oɇ*�y�A)	@��Ꝃ�˖j],�,���Q�]�G��M�alkx��C�F8.�Ge�!�Х�h*�.���{��7EŐ��"@:��j|:��u�.@FN�C��k�=�ɫ�����!��ˊUa�9�y�Z�p�mӥV�uhb����͏.��Mx�<�ģBq��}���Z�������%�d�$��ԉ�4�%�7ϛ7���/������m}���9y�����Q�YSJ,������M���(ȹ*T,b�>X+~9�Eߝ�x�]fn��Գ��a��x����jnQqD�聬�H0�wѤ�d��.NEk���<�Z������$ny (� �if���	���X|�{Y�5ďܖ�Wv�;09/d���@W�c��;X�<H͓e<J���K���J��n��[u�W�i��/��n��0�h���C�ߞ�^���63l�����N�~]��[O�Ml������ڬ)j�G#����J��)[�\���Ͼ�}54�Y$旕�w���&��;{(�U;yJVG�W<jdV�XR_��SЬ�!�0��k����݆GU�>s0�Q���b!2�{�8�X�hCL���;<E鯽,7�a5>���|�xܤX�!F���e2�]�)J�A/��<9��Ռ4���`򊠒~��������˜O^;���}���J/AA	#������Z"L>�������>��/���"%,bȖL��ծC�vc��!;��?��!����$ZJ�`Z������yM�k������ٺ߫D�R@D��N��V���8��p¡^X�$	P�<X_�����u0��6�+��#H��s�˂T)�kvd'�98i�VA|�>�8]�2P��0Y�~����Z�t�q#v�ꤷ���J�Yl�AG]|���IV7�4�_>Y�oCN�8S�6@���/���D��ߡٴB�)#e����8j�����b���<��k�$^h���^���d�M�~�A��|��}J	;������yp�{&��U*��z��^M�f|�����?�3�&�h�$��6u���k�jJZ �H�#�I�/a����~@������-�V|Ĝ:��:T�]�m��(�6�ab��귢1��mrK8����̨��ǻ�\��G��Q�a\]���ΐ��"������L��'��kA�n�����}�KhPf���֑����'�DV^�7��޼�:��{"�)�\ABi��KjY��� �1�p������I���22U��RX��IZQ��Ƀ����kڪ�nr#�f
�mUgL]:&].������ke�gs߬���K��p� ����@���O̷Q���v#��ťߤ�z�ه����E�sF���}��E�5���6e �=��Ƈ,J|�٧
�"m�vT�"i�f�b���Y��bس����5��#Iq"F[���P �|Y��3Y��}e�J5�`.(-3��L��w���}
J!ᨮ7�>%���`/R����L,���*�@��nGAP�@�7(�Q������Q�G͢7����I!NC����9�]L;��pf�2uP�l�n�^�����U!'O{0�g�)*���-��u��Bs5���&���Z�A�H�b�
�a*?cA#��Ԥ�����J	���x<�I.� ]���c���5�e���1�8π���v��[ �J~���M��I���~j!���҅|siO��V(m ����)5��e8�G�kX>�a�5�_8t�ջ�oӗr��sq�6��6k��Q��-�P�U��P6(Ţ�p�]�˲���7����&HV�L.N^�:���g:Ĕ��Nb�KI_��mI�׉ �6��4�����S��z&�oe:?�b�_���(�H�MQ(41��Z�b�� ~q-]#D�Z�F�/���6=���p��"�	�v�W=����:e�QyC�}��U,R����{�;u��G�N���I9����!�P=��i:���Wԩ��Ღ�5m�:�A��_'n�
H}��M�>A��!��x�����%)�^t|7⢰-���?���ʦ��ps��2������S&��K�$R���.�y�����$|���FX����}+�*�T�*U�qJ��!<��1�R���Jل-V���:�zo*�=oo���Gbr���A�]�d#D	�����&���Le�f䶡�������ؚ�VS81Ѵ0	��O't���%P�h�Q��><�b�ָ;i��]GW��e7���'эȝU����f��84k��q�d��ER��OC]j�l��H���1[@���J1�ZY)oM=��n!Hs:x��/��K�j�h�]�
��,\J���Y��|�w]y��S��_����hq���"�({�{H���1�����fu���uJz���ʝ�����B�_:��L�2��wGH׶�.�a�0n
n)u��z�`�4Ej�J�bD!���G�p`���VA�#�����^s���} �z�$9����2�2�
�X��Rkk��	8�>]��l��+�;ޡ�.!����5Z����!t潳}v����m��^z��κ��x<Dr4�ìȞ?鎾���O��g��51����N����?,���S���!�R)fd�����+��!��r�H�Joɔ�w뻢�	y���S UT5�c;����l=��&����4#7Q��l����dl��i�
r����b�t�͑��82����9_'��׃��&#i߾���V��0�䜐�\���l��ٵ�����(s@�i�c�Ǟkj��� 
�:��̊j��م@����q�J떫I#@di�	���{S%p�G�LZ�hړ	��c�%M�\,^��_9
��W��n�nT�~ 8?x���!6�Ýj�כn� �-���
��5����B�p���L&1�M�cT�����]�������6Ȳ`퀎�דg�%x�yߐ��#t��q��6<��B'ZM}֫�AT믺?���;��1�ԹLD��_E��A1���F������|�C�"p ais]�K�g!��K�N�_GJ<v�S���	E�.%�:���N���vXK&7�c䳽e7�Vs�s�Il{3�ԥ���|}���+L	Ą Jq'(��_��o�A�$ 3���d̰Xݝ���y$Y����[��w�ɽ�%�)�pT�����>�+Kl۪��0�~��Fگ+i��c��o�c0B

I�����w~t �l��~ �a���ylM)����i�K&�~]�£|� �&�r (�fl$���U���Ң]$"	ـ��-�HJ(�'0��~�lCP���E�'���O�z0N�l��$��NUv����D�K�2(b�ʌF(���+�|�:(�R�"��|��\R���9ܸ�&w�#g}ÓG-��h�ֵC�:fp�j��o���A�p�e$pI�z3��-��-g�-�{� D|3�ݍ|@�E��������#���L��Z/zGer�n������ç�p��(�p�kP��Ú3�;�酁�T(��-],�k��mۄlE�j�}�@�׶v���wC&MX�b�N	����/i&D���'��$���	�5��6�L����J����rY�����Cq<{Nlꗇi�Wlх7�jp�*o�Q4N�ݺ�8Nw�&�V�A��O`˰�9���:Y�+}��Ǻ	�c]�ǫr��+�"��`02����C��dV�Wf�Rs��f���^�ZCq�c��D�k��c��B���V?m�;�xy�˿��d�>ӤEBAP�/b��k�z4�b��lG���^m��z�3�r\�;���\s����=���MK���	O��������E@����S��f�ˠ]�FE}!�݄���igF����an��Z����W��c�A�}���������J�v�����|�x�%A�D�b>p�/��?v��x�����1��o]q�ֆDf�b?VAd��D�bp��L	wsǷ�|���p#���DPhB��	�F��#8�˃�8��i���a����P���0�li��}Iq15���m�sV�1�C��>י�}5b��lj̻J��A�.�)�&%{��qgN|pa�ΗS��֔dc�ǡl��;�sA��j����Y�jš���&P�&z�*c-t�UxU�w���Top{PTb뱈��X
�t?ϐ�5e��QXDxi�c9!&U����~|�����xKtc�V��1��ViQ��8�[����0��I�����#z�����t�VF�������;[��g��LkΡ���쎝�j��ˀ#�H��丝�X �uK3���rv���g�I	Gj�5S��1��3�\Eח�S򣌅�COGuS�޴O��a���
���@��S�}ב�o}�e4��϶�A���7��_�k��T84�R4�Ѯh���Ҧ%���&��H˙M�Ÿ��0��mm��s��҅�?�|��/mv/�{�B��r�G
0ucpc����6���:�Q�SN��R~�	Zd@���e��`Q�����w2�l�x�Ҡ�mٵ�^T�~�VE��-��=�����}�u��p�,��l�B�A7�K��|�]b��˫���t��s�����jMׄ?�Ի�Rk呴w����O�Y{�)��B\�=bTXR8���s:u�?I&m�_a��4uKeZ�g�W ��>��{z���SS�!�]��^I�J�N:��#`]jtj�@�c��ɌV�"�Q�BLS��Z���}�c�~u�UÿN��^=T�52�y��S���d�|�2��*H&�q��N��ޥa�Ul���-n�����Rݫ\p� }�pIp�B����Qe��4�MB6��h;�L�р�JM���?�:B�|�Y�^kDG�Q�nˀW�lq�r�|�?맷"���T=�|�@9Em�*t/|��^ku�
�s��k_�)rY�t.u�1���#�qr+��������F���>�tik&�z�dM�H���Dŵ5����Jk:�X���t����-ٜ�}RL������\�C>��l�;q�s�v�S�Ųh�������-�;~�g>��ɕG+�W�K�[�r˿��� �s�`��t�Ĉ�ҁ����7Eۥ��4Z\dj����w�\���|7��"���<��l�>j������M�O�S	�����G�ݠ� �]���D� w:Y�^T�H��"���*��|��D���Q��,��d���1L�^ޜ����{�e-i�f
7����6�B�z���u�����!Qs��|ˏs֎�c ��󞸜瘭��T��ކ�j�a>��};��@�4��PW��i��Eq
zd�j�ǭh���b;���n�<��T/�ʾ�<��JF�.ŗP3��wJ�I$���̓��l�E��cd.��d�1�y��V��� ̐�eS#ÊI>[9'���I���'KU���G��4@�mz$�$�����~M(�G�cm)��.����pBD��1���YQ
�²�"��9�'��>��b�J�V_n��кc�Y�+�90��?��6h#@�I3��G������m�Ń� ���Ҡ6����>�'���~1g�����4��`���'j�VoS4�N0;�]H��cG-\j�|�)�?W�E�Y��_`�I6:��z��xA-DP�[�
�V�ʈ���e�-^��-��;N�����08]}t�*�1�S�Q!?��X��,6I�K����md�`�_V�~֧�����p�﷒�{�J��R2��j+ �/]:U�� wnC��XC���2/ѥ�2E+d�wV����yzkQԤ�}�v} �k��4l��mZ��� z�PO�3��Lϥ��Y�Ν�B{��g�&f���B'�3f/���8�Sj��[��I�%�nV��ݮ�R}a;�:�Bz�%�t�z$�6W��2�7�i��-L�t�֚c-Pڧ�symܳ�cKKH�"���R��2i �_2_or��y&hn+'A�˃W���V+�;��l���
�al[u��@J?��
�ĭ���'�)��[(a���]\O��f�pz�=��0�7�8l��R�<�gjF
t�A��ּ�%�������r�CU3�虚�e�G��'��"gC���c�W��M#F�y����`{�8(�P\(U��B�����f$$K5>h��lo�c<;�1��t��X�K{�"��r"�8��.�9i:<��k�XT.�%�H�b�SK���b�!���2[������mO��!���4M��ivBC$���/�<����4i˟�a~/�	�"iٴ-a�+h>	o�f_�T�ꭽZ��@|�F�fx�]1}M���Z���M�tA%5���Gf�el�|l�N�C�Ň&�$Vb��ó�{�oo�V�t�-r��<t`�"�L\���,a[{�P���Ai�:��߯����.��cf�F)�쇣�S_�qh��#:��b��k������EfZ�*�B<�a�> ���Ã�.�`&~S�ށGX��^p	/e�cV#-��:K��fQ"Ү���,&�#C1@ԚZ{}��$�)z&���@�J&k=ч��䌋�j��7q�a;t��C3�Du!�䷺��
G�W�?9?��#��Yƭe�`���'@�nm�$�a�
�ȳ�0�ᕿ��F�����"eb�{�*+>m��y�x���,ﮪ��[����7��XU��A��aט�"flq�J�\�U.)�W�y���C;s��,�,��w@��n2<?}jO��3\9��Bv*�EK�������͒����tl����I�ǥs�4�ǎw���j�_K�.'�F��5y���Nti�w�:��q��[U����'��P*����iv�+�;-�O�h�lj�ƕ���Ta��������z��-��d�NPZG6L'�g�c$E6���r6�e��r�=n	:8)?Я@�s&C�ԜB�IK��)�3��ȥis�^CU���#��ֻ�$�n?�)���`JR=��H����÷ҝ�1q]��?��M(�-�-]$e�a��.bi�Ó.�j�T����FxFd<��j��t��~�W��N��q�L�h���%9M�S�9qu��[���W��Dh�ͺh�`"^Em��U����}&��6�����ڄ���%��WF�U��f3�B<�	�7���H/�ð�E �􆿃�JR�O��3�����g���\��6�S��l�Y�MS�LY�S�)�{�I�!�cʳ�!I��t�F��%Ԝ�2��ST�G����e�w(�j%��3�H�U)�Ѽܦ_sFm�E>���XB�Ϧ�67�o��ʹy���eV�����)���(�9MA"Wg��#'.]N��&�@��5����:�8��g
ぽBH{�(�;�����Ya��
�HS����3@��R�r��ă]�`����y)M!�{t"��
$�$�5��*�<���)�ᐛل��f1�ad��@H�5������h��
C�lP9�>��@�v�@t9�G��>�r;\��)����y�B��%�
~7\�tk�~����S]��v��N����AKjH��M��/U##:��LxВ=�Y�[���y�/�G�asj*^����ގf�i �h��fRj�����7/ ��[�I.M�cC��1�4Ĵ�&��f����$'O��=T��`r��t���\��t�d��<�+�яӽ�Wk����kMın�?4�������O��B+N��*_a�(�'�rl��pY,`�.���%@o�G��;���LR��qa�R�K�3��=EW-M�u�2%�z�B�[��>��c�����dg-��=T`��j8۪�\>���.[�Pb^J.��ԊoT$g==��������e��(��E{�x\��^Q�Uo�}u+�y3X�����u�}�\Pq"�B�F���v�"ԋ�[�ʠ�d�ǐq�Y����E�°��֛_mX�(3����Ej�|�Î�Р�Ή4�����eؔ,�+�t���W�Jl��'��0�X�h?e��I�l9	ܚ$�Ci���1Ц�=�Z�9/�!�\���<�Pp~�c�g� ���i�ޑd�{�`>�b��njR�"T
V�%D-*9���a�u��IT.ŉ����I
���`6��N�CJ��CMw�ߧN�^G�Z�+O3L���Ou�*y7��~�"9���gq�/��{�@+I�"P�L��L���.�V1�An���G���"���`"�D=Ss�A�re�k�tY\���2{��+��;څP�U+pޖ��c��a�\�tO�~{���U��`6$�12j����EJ{]η�jB>|��j�b)�0F�0��@��ނ@�)$����~DC�KU$��@♖<��s7��`�.�0���֡��$'����;����B|�]��r��EFg
%�Z�j���-挅���,EJ�-y\I�F��N��'=�H� �S�O��C�E2
�]����!L�73\)ο�K֧��x	���&�I^@6= ���MkΑ@I����ds�`��mlɯ��w�([�PS�5t�1��|<�O��FS�6��1�f����_F��=
����u�n���\����ʢF�}����.֚{u����������s���,X����|��n"91��~S�I��_,h&�28�|�|���če"�n�]��_��LijK�ZqӺ�}	�,w�H^H��v�����W���J��7�)M�AR�]������|P4
�ҏ� ���>#�1�zE� c�&uИ��1J��$kP5�_�/:8���������à�y��� �RL�7�\���)�����	cFV"�e��n�����]M����k���Q���K��>�2e�I�ors��UGzf�zNą`y�L}0����B@Y�.S|�G��Pi�<����A���}��պ�������}�[f@��oP�*XMb(��ۈ�V�U�D�8���(�P/��Ft�b5�l�����r�#?�(\كM��lMb�����^�8}�Ny�	�si]	;��a�� �q~\֤�w��8K%9�촕\AE�@`�^��_׳�]���^������Y���\Z���-��2���kj�uD�		�E��VK�?�s�|�������g����gE�v��:4�Ć$��䨳Hs���Z"�Q��߂�#��մWشjZ$�A?$@t�K�ĖƢ\W�d����s��i����,�J ��C7H�>D���e�I�v�I�Z���l?�t�<8v�I0�%|N�E>�;�f|�Ŏ$Z>,#�Հ��W�Ԭ��D<n&Ƃ�9Ve��겎��pCǯq��$��"�t?lӾ_+�����t'����m�A?�����HƜ���9;/��Ո�����E��<m/zs/�b��o !˹�4W>N,iY~�o�)���z�\L��(L~r
�s���X�s�˪o�m���r�"�?G�Z�$k�ѐ�R7��\����!�����u�#֪}�fTBm�c>��@o>'g��w�O_�.b�q\�+��9�lM�4RyCY�H����֜��U\S7�����Ϸ�'�"gY��)�:�j�~9Z���Z'z:��&��Tl�m=*f��m���"!��ȵ��z�?�Lvx1^	;h�h��Q2����j���1@y�Bf�=�=O�\Y�*�~a6c��m���x<��4�W�g���d����v��Z�\c!CU�H����L_i��;ھ492?� U7h�*;��Ƌ6���>B̞mHA�b�|�~�U��'7��ޛܳ�*��'���&�է1�{���Nt�t�C|FF��;&������!�����R2T!���V���l��u��D\pV����}���&��`^É���Z�O'yϧ9���3�lke!��z��(���Әm|��-�.�������F��c�=���u����&��b92D��9��^ y�����@���~]'�@ y\�4�T���&�u2zp�*�6�W��U�FJ�}�9垴�2)�L�T�]u(KD���� H5�5I���S(j���9�#^�%�~T�^v��OI�^N.Z�Ǆ�x�N����,���jSa."d�A�/�a�Y�18���W���;���V���x����(��Z�s,�&H
��חA�w�G����B��8�~�&78�,�I܅���S�����^)����عM�[Q�`��ɘ�l)@�g1��8*��榲
��*��C�gr�����c�vu5�,y-Ni�.$��������Ĳ�k��S"$�����iu�+�R�K��٠4���!}G�Z\�T/��`���J�R��qo��(N߷�gP$0�!�/F��K��	�L)w�P�N�$�L���\l4-���3�U�Qx�|�\2�<�@���Z^J�>}4�*�I�h�}4]D,v����o.8�X��~�n���qyB/�x����)�������Nq9=o2���������*�>�X��f_{�,���odaO�����
�w�~;��ll�T�S���C����[�^�m���T�^�������A5MAz�>�_���S����1�dv~��c�@��m7�7�^{�?�"�K��8k���i�1�"����[&��>���Z�����ʮ�j�?�E�v����_�<<��0�m9m����-W���x۷D��⫗��G�/s~P�SF47��'6�}�K��Y�Ǻ7�������Zg9�øF6C���� �Sk�F�z��Od���=p��fzd�pÃ���0�9�2�
�� +�b�G�Ke�!ج�T7��G] /@��YJ���$4_5� �\�u_���� !�R�k�,�M{b�n>�$�j�Z�w{��=��c��k�-?2i�]�1+�*H1��y��mDb̘!��'~-�+��������b�AS�%KA'L&�M�I �[흽k�;D{��/�&�]?��'$�D��Y(K&��M�&o���':�[%�iF_֛xɊ�=�D�f�ǧ@WDN�]�G���j{�}�[�)B/���	"���U
���������	�J����� �c�Rd� ǔ4:�N�a˴���O�rxoƦ��M��}�N�����Ď�@X��z���\���z�ˈ�4��,����ݡ{����w��H&�r�L	6�$���tV�w5� ��=�u|��w,��͏�գz���F���~�����N�	7;�!��p��*go����g]F�#;u�B�������f��0� ����ҹ�{��t~�d���I:K#�֏�Րڻ�ϠB8��:P)��s��C�ӧ��F�+��ďo�-1�����6À
$�3�=�%�wЂ��Z*Q;ަ�l,;�_VS%@�G���s���\�s�S�ܼZ�n䔡d��#읕��s[)ְ2=�"���|�`��^�������TbN�ee�"[$�y��c�c�j�Xǐ�@w����j�8 G�QT�;w���c� @�+G7:���X�"͋!M'�f2��Nu��t�`{���Rw&j�\ʮ��|౥t�[�y�Y�#B.�/l���<��5���CG��������O;�Z�ߜ>#P��$T���X�}UZS(��r	/���N�աgjCiֳh���>�'�*�{�vf��+�jo�V��+���ͮ���~�?��\�� :ꚮp>��{�+��|�xO����|��S5)ȧ�	U�uT� k�I0y+�����f�ܶ�W��1Z�=�C�h�K��/8�)9|g�_�	�lGUB��ܛl��sc,a�(m=�up��q��DJ�%�S�~>ȳL��0�bE�Κ̹���D&N���:puho`�g�����O-���F��m)��o[މCo����h}�
�W�����`_�	�b���`��r��!�ojSn%"�z�k��)�9�e5����9�Z�j�ﲵW5�5xk+�q�֏�2������<"�yr��7ek�p#�cw��=Ao�D��Sk1 �P6r�/�oK��}qmӤ�v�vt��^�8���zM�*Ax�&�5"'	@�z֏�'q�(ܛ��'Сe+ymL�-��p{R����o�R�C���f�c�h�Mƅ�23_]�ƽ������1m@U���i�ǯ���S\��"}����͞�*u��P�M��q��Aq¶/�T���.��M��1�(��^v��赀aD������Չ/�+f󨄺X���o�pE��t	���AT�S�ޤ�s�
>$df�4<�t�s����Qm2���a:�e"ʷ=jq��^���&�	���[45�!�$�"�}����M�'��*�y����KTѺ��m�j��8bb�kZ�L�?���M�ߏ�c>o��+��!5M>֫Z���%p�fAEQ_(�=@�xo%�0�ha�3�	�ic(�J��D�P�ݓZ&|�5��3a�&�>��Ƽ��l����;z�ΎK"2)��a~�t}΄�nuL�b����p�"#G }^�X��U��5�����!�.�n���8������~�d��(��~!Ə�q�¡1���͟v��Bg�Q���� �f%����?����த����3�J,��I��)X��Rķ쮼J&��n��o&��\?�\�+w��\�34�w9,����Q��,"v���X}�]<���7d��D����=�}��w��V=�%<��T��d��W�/�/O'TP}w��h'�i��b����#�![����AX/�z���t��m\S�%�0L� �����ǉf�l�X�)2��6��*���b$h�aB� �{Чe�
tfF�.T��r����a*Ě��]�?�>"���)��)��6F!���AzRtQC]~���Z�rJ��_lک��h��c�oO�2f���W[- v��|�TZC|�8y�;��.G��|�ܘ�z�K7B�8��@�OsJ)+[ڝH�ZTS�
�~���Vܮ0U%���b�Zr<���r����h��b�w�{9|���{�h������ހ�-���f4N�wHۛ�� 4	,�ڐ��"���HB4��>�-?@� �R=�="�����(�~����h^ܳܬ�r>',���T����1�4�*R?��|�O���*M�
@Vu��|\o�
�Yjk��;-�E�� �SF3w��4�#�E]؋����2�� 9m)��B�H��~ qVtG�JT�!NmBjS��;-%xI#�e�al��Ki������=7a�w��/�5�V�<��~{����L�����O�kV�QF[ڐ����t�4��X�����Y��NVݯۭ����Әhԯ�/��^����nA��G�)_>_�;kTQ�gU��� �Q(�:Ҋ����fn0=���l�e�SRH)�t�њ�ٍkW3�8��0eF�1�M����������	��k4N�����>��-SK5��@���g�*��>��r������iА?�P/���R�(H�5�y`�q?�*>�U��1��n�Ov#�Ӊ��yn�D��p��|S�]����Vq�'��C� B��������F����o�}���;����}b^La��|t���5��������Dgd�X8�}\���rnyN�P4c�K.~��
������q�jҦK
m�QO��ͽƹZ�@�.�<9;��U�@5Eg#)���w*�;+<����M��GfN�S��6D����I;m�c����<.�i��20�	���RtC�@�o�V�ڝ��D�?���R�R!���
�p�}Q1�3�$s�-�g�?�M�m��r�ur�6�S$oW���)�T �����xa��53D�;c�:���׺��<�_�y�����nÓz |6ì�
%s;�7���}�;��[��<�S|��k4�Q�i5��*7#���{ǃo�`���橠�8O<���zM�I$@ͤ�aa!�^M`��5�S[<q~�:2xl 2ͽl�7/�-�F�����/� ɬ��:o|�;��3G:�)�䎳\�e�@ue�:�Δ6���钗���EWZ w��<��ڳSY�a��$>���L�H���e�ͬq21����v�� ��a��tU��b�tJ:�������"�fF;�Zȝƃ��Z��͇����eLk79Z�?I�w����I7Q�9�+߼iOu:�L���6�0���Rv��3в�k��XDY0")]��S(~��� V9\���������j�[���.6���	RM���:���5�"/QٚcF,K��!q�#6���i�ψcy���@�Q?T����=�#Y�wA��r�1U?�p�5=�i���3*r��U�1��,���N:+�6O^H��ּ��o�O\�:�t�S6l�AK��nf��/��nr/�kP�&�"��u�V˖ٓ��A9^qr�T2�� ���٭�������n�P�g@�[M���l�xy+W��%,W8_%s�*�����r�&�A�_k�b�9���4���C����W�ۧ��9�p�����4!�`=&����*$�ܡ�7�l���%�|��*F���R%�w���<K��K9<W�� Cp�b���!�^��xeLx�kw<��(��A��y����Tcɣ�ª�a�7��g����5gMR"�yIgI�Gl*��+R)�qu:Ym�����$�>�>|n��-sL��Ɯ�ё��i�92P��~ke:��ܳ�L#�d����rG�G����u!��	TE�H�$w%���	�w�P��_���!��H�P�"E��'s����:��d�F&٢�_o�C���#ˀ��Օ���ivaⅭ�4�f�alF�P� B�VZX�h��ڞ�\���#�'�K|�ib����<d�vI�ٲ�Ar�v*تT��ox�}�T4�5��ķ�ҁ\��i� �yT@��������G
$s��tBo�X����v�E�Ո�QQ�z%��_�z�G(_�5����Ke���E"y���:�\�d[�sV�����HF��)L|����xlP�L��������H���-��o���2�\-.�xA�^-p
 ~iFI�h���%m,�a��H%��g5fM���p�<M��e#X
]?��Y�r�Hm�-"+E��oġ��3("��1+$n��ψ^}U�c�w�������A�2�m�>'�����H�JJⷃ�I������#J¶u�@XC2K��n��,%[?�iu�u�=5�c�>�T�3~��vf\����YYԠ.oyx}�;"&�[`�M�i��ε�H+;h|�������kq�_Pz��8��r����m�J�W��1���m������/f"��J�r:��8Ol�E�b�S�E��[���|N+�(��6wZ&8(�niE�4�^�I6B+<��?��eN��-�ُ3��8���!x��~e��9�Z���P�B����]���\�;E���@��4M�S_L�����|a��6�F��5?����~�h��\����q�d��@k)�~^�!�a�ޑ�\�;תּ�^��]E)��~�@�v�¦pzK|-R�K�Z�߮
^i��r�Y�0	/B�وW����� �e	�.�Eb+E.�c�9��{i8��gjf'L��=�Ԧ��?���(c�eHV��kM,�[@����]E�%^ Z'u�&�;b6�c�I��;�|�@����l�=�v�,'�Cb��3�{m�_�I3.�ʼ	�21T�\(7i�����c/��m�F��
A����� �I="k`�1���c�	�����3�'�1�%k:�3V1 �}Ü#�������0���� c� ���Rr�+�r-�`����5�}@�g}�)(I��="xs�ǈ
��|�o������V@���I��Zc��#��n�(��V5�_�P�>�,sL�<��\^���uV�O�l�f˔�v��cqڄ�߄�S�4�w��UD ���7�O[�<�2��bJf=b�F� ���_x�����D�$����IT&ך �V��EnߪPZ��L>�%� (HH�#
M?��]���8��̓��\�z�_[�7\;���3����}ys~m��%T��K�LD��4�yo*k�\@:�0�6�iI?����ۏ<�c��5��X� �˞QTH\���
*��u���e�}���IdW���5�>�J��۵ʾ8;B��$��v��D�<����y%���Z3�.^��.|�|�D
)�ǻ�I�]�e/�f?�;��$u�2̈́��N���K'<�/+o�����;*�xD�NyU�7q����y��, �ߓǆ�K�����hfx�ľQ����b'Xt�"�wM�
�ǵir��/�R��M�2G��=��H=�Y�d�"l�~�%�VD���O[�'%J� Pe�Cgβ�x�'��Ny4�-�6T�<v�LM�q��h���A�H!>R^2�@�l�����;.��/Z鎟҃�� ���H�X�EO���G+��c�cVUQ��D��u�'b	�3\�T;��
�#�9�:œ�5��>�-��F QRF7u�Β��,�}��)��I��yT6G���q�ֽ�4�#���i�w�X����>����`�oh��rru��y?����M���\\qr��(M�\ބ�-�qq�U2w.�b :�viP\�{|�\�g�]?t��5 I����摔w�CO�2��~(g8Bd۸d�s��&,�D媂�w�(JO�`���^���3�NJ�)�(B*�㠍n���r)������ώ�{�6�
�0֌�Q�?:_rJ�A�&��9�=�H��X`���&* Nl�8��ؖ&g%V��Jzծ}n�c���q�/~ӓ4��Y�޿+?��/*��ע����)��D�����h�mY��&��o�b0��-����[�4�h]�5-�y�r�0��7�K6�{7�������sC�Z�31�u�DY6�?��Ùì_����m�e��r��
�n(�k*zF��5���<����B��C��K�:]�{������*�7)�P�!��k(ڳ�8o�3M�q�/C���ӱ�����w5�̟�}���Sj׼F������-���1,`ѹ����8k�;��NDZ��fE�����R[5}w=�_a�Zln�z�`���E�Y��4�d�Њ��W�H�-����Ǽ����'*ef�[���gM��|��)���C4����f��Z��� jۧ�D��M�2������ºP�	���@�>�_�C��h����5����L�LÂ�(��r�t�k#-����{��\TT^�U/�孪3:���v�p��C���(^��č���5��o)��:_5�橜5 N�5֍�(�G#hd���Ţs�'�V��'��g*A�A��}�1e��l�p���V/˽� WKE�(���dl�L�~;���M㤍��9�fWN-|�d��n2���zҖ�I�q�L����P�i�ѧ#c�4�O�(��rEH%�<�hQ���ۤ^�d�pn��Lfu�i��<}�N�|K��哈�_pZ�fh19+�� ��iC�xd���5��y�^�jzEW3�Cq���]xn�HVq���Q+U����o�$I�t�=�w�~�ӌ���O��F��X���?��)ٝ���"�������Dfb�wc���2�~J$�z���b�"� fa�m�\�co�\����jt�Yl	��l��=܉;��^���PL��ޖ�����ܩ�Y"hu_�^�ws�!m{�o1�8�a1�����|��d��A��u=���Ǩ� �5 F��}�S��op��-�f>l�q�Z���ZP�!��F��Z���޴�7l+D��`_�ZDA���
P��i!���iIWn�r�%�Y���Z���b���������<9��:2e���N/2�?�&���d�sg��[�q�(f7��]�1�&�>z���k)�EL�ͱ(��8�p�?��{��A�	gxC[�;w����}Zԧ� �TU���6"��W�+U��Y�;�����1�^�KFA	K�6�u�gݕs�eĄi�A��u�h�PH˪�J�h��X�JNļ_�N��'���N[|w�]7,w�J��+'h�îxX�K}`�CWr�bc@� :i���f5܊�9e�����M��L���$F�F_��MY�{�7ٟi�����]Ptns1��P$������\�YWR��l��f­�c������pẞSUzSs[����H7�����q��,ouAB��aFw<��bP�q�p��9�24 ��?�����!	����@R�=_�θo�h�_�I�""�H��
9���~�ݛ�+iS�{?8g���ȗ��!�VZh>xԻ_���B�ٮ����L&���	��PU�M��ka�ͩ��L����go׈-����X�س�"��e�-P�j��j�\<,f�	2u�'L�"����>�:�ƿ�9�Qz� u��Hg�=�:>��N55`����2�}�VD��m�Cԅќ�;O��u�N|�^�C.5��$L�1���@��$+ś�"z�Z�F=��c7�ԛ���*x����].�@@�X/?c�;����G����K�\<�UAo�ϐj;]bo8v�Ofg��r�+�3�YD���3�H(�1S�qL��C��5��Q#5�Fڐ���2Ku%�������U��F�E���;,W' ey�Fg�w�d34����8i3��b0A\���`���{'VzD��E�&L�'����艬iӦFw�����$@��Cp�mt��5�7f�T�d��zlAdu��L�1/DAdO�,&mU�:e���� �M�UUU`W腣��(L�5-E��T���
[�����3e/�$3�W�����H���p����1�G$��Q��8��u�h"�NKha9�/���� �p?2Q�̭>����R�*���q��r5QӮXQG;�� ��^S|i�{�Rd�p+x�XT.�0�s�)1>"8����fu�Ht�C����"χ*s��)Zj�4:�;���u�xNҔl�	�~[C_+<d�T�3C9D�<�d_j��7x�jB���_�oݸ)[���CIPQ2ߤ;�k��$�{���㿴�6�� 7q	��A�=O�|ӼӲ�����*.h� ^.؝���db�ZZ��ȧ��YŶ~��&*,v@�HKY���5'�N�a5���n�|���.d�-Ls���]H|C� v{��7 �[%��_�^�M��TAth�\�:(P�Cw�������{/1)W�+L�����y!�dU@O�Zt7���Ȯ�i�g�,����rY��fXca����p�#��畩I�W؝�q�<ؠ~ic(Z�P$�!ϺF����*��Em�	�K�Á�Ńz�%����WukѦR��r�o
C��߶	��P�t9��,Ɛ��5n�
����+�m�'�S�!������V���
<}��P�����n/3�:E[��	,q��M���K���ޠ3!�g+)�W�Ul�o�B5�w��hK���%�u�F��ڃ���B�����Np7�X��E�h�{ь'��bfs����&!x(�l���5�v����3��ゖ��q̇f�$4�M���5F.�.@L��a�����[�0��Q����"?�&����u��m�R=���4~�CJ�����N)���I�j!��@��N���f	?t�MSz2H�-�xڞ�`��Ť�P6�rԜ�؏9�9�n6��x�}��<scm�Д��:���9���m����@�3�����x��v1��N������Tv�|��>^8�X�&��mE���K�k8~����)�4�&� `��|9�e�zY��m�x� �����b������b���n� ��ǝ�jf�Gv/1Lq�ĴM�Al�ǲ��t�K<gS�j�j��XK���4�(�cHzc�cL��*����Y*�ʊ��,/9�4'����Z��n�}�l�Ӆ�t��?rg��c9U�`,�n	����p�O�{�Eߟ$�ʆ }�D�j�bU��h#>�z�G&Q�m�{a�qL��>���S�Ȕ��G�1pU�\�?\���G���!�OPJ�lV��px����:S�"�AU��A�B_u�;P�*ƹ."�H߈U��B�>���d��]*�x�;�7"l���O9���iPv4��9:0FK�����^�kH�"	{_"�б�u4n�34��*���Z�N�����>F����r�����9rf�'���?.8�$�
� �xc�鬨�ʵ���"_��s��Rh�:omv�p�%&F�P"ǩ�\&�U��!oG�A�����_��P��ÈC_���Ca���u�c�?�� l�.^q��-�jE���{���������M7`�Mש����Is��qOw}��t�&�+���P�*_I!ή�:�r�>���쁩?_	�M�W���zr�Im��y���Wc� �^+`�q�~$η���	.��?j%�h��׈N��8M�׶7�d�܋e�U��v~���4�x�i��OA��,�xR�g�S_�<�I�d��u,�V���ÅcS=�PB6b0H~oU���nF�G�>'�R�#&���i�˂��5ի&�_��\��P�I>��Y����[0!<���y<K>���5��<)�� BB;7-+��{��b�렍Eզ��d��Uw:_�1�'n?��5� q/\����}�����2��k(���}�����&y�rz͙7�9�w���H����Z ��<��<7>�WQ��?*R��W��VK;���7k�t��4���K ��=��3��$�h�O�r�K�Ɇʼ0q۔�f���#�,e>d�:��3;��yթ�Xq��c0es��o��A�Y��!�����/�ͅpp�3�m#s�2�f)8�~1D@��%b�A����_�ۣ��XC�6 ,��]�į(4	��@�,��'�%
�:'�5�G��Wt�wm�R{x�m��]��]�-i�T��l�!gK���~���r8:#��]�~��Q��<�/�i�Ѷr�Q�m��R�C�w���Rz�LäC��@����\lo�{}}�Gy���'8#Vv�����4V�L�q�v?F�x}�{V���Қ~�Y8�z��m��c�>�_O�����N%f�X:���O��d�$_!��T*��k�/�"�8&��Ok��k=Z �2�W[�ZWb�y 挻�9�[
f�"%@K���9k���=�¬"���l�h��NZ��.��>�ނ�yg�ɷÀ���+����r�0Y�nu)�+�'��W�4q�^X�H��5ij� {�hnU��,�ty?Dr#S ��D!�G]0@�P!��)FR�|�=�Y�, D��|vB�s+�%9�<D�; ߷y)�7�h�33y��0���`�+Gp�ec���$_�
ݘ�/��a�-��tM�B�<���B(���dҖ�rv��`�ƱY����p������k��k)�d:*-�1�8AAFD����va���A�o�z&�F#��?^��D�S����'d��R,��1V)x�I��!��d8jPO	�ɪN�34�ǈ=R]_�>�dflI1�'>�l���BbK4:��\�lj�e�Q���b����7-�&�^�i���ؗڛ��ب����1�Y%9ht���PV��_]3m��\�y;ɯS���PI���&ɤ��d��,G��֬���>������h��`��lI��ȅ,"[��"�>� ��r�%I�����H?
�AY�@�%�j���M�bi�5��/b��q��U&�}�^����>-���"sib~��*�4m���!�,��->��^0��l/tO����n���	�G�yiq�l����NB4�9�B�f��Od���M���(:�?�.'�oߎ���$k��E��t�ڦ1�Z�]�h��r���D�Wi:Bx����&1]Hl;�'-�kK�_��tL���8D�\{����T3{0.a�uWZZ�����gl׀7%�Pϔ��B��p�#�W��7��,~s�Y�*�	�M ��;��MQ��h��rO#}��1v��~�¯!i��\h�� :N�QR��T��J�P,w�ͽ���!)�0��s
��*ET!��Ve�g�s���C���ߐ"
��B�F@�w1�DG��i������A�2���,�az�?3<�zo$k�*L�|�Č�c�^�e���b�E�{	�U\|$-�N�J���'�FBK7�m���`�\�:���R�G�8�#����E��8����-�`���?j�'�m#-o���qX�l�S+���m?�ȵ�#�BF�+f�lR�C'̊�MZUfX*3��AZV���5^0=Q��<M%0���� >�Z�d�\L��l��d�޽� j8ĩv6W�i���`o���G>b����Z��0f�K~��='5 4l�j.��e��N��#-JHn�P�~��?�o&r���	S�Rm�;j]��,��ܲ��i�!����k[�ӎܔ�!�W�ʶb�>���&k��JU(T�V��/�j�P�/C ҉�!�F=��p�f�7�����#�Y����1kz�h�$;ok�i�ށ��'�qO�hr����b�*�ST]��H��W����x��|m�2������JU^G�����Q��V)������/?W��b��)Ή����M��s_����X�	v�J�(�I��T��Y��:�J�(Y<�g���+J۟?�nJ��sEq"&�'��i�8f�n݂:��YR��
{R�l=�nw�oE۴����e�I��t�g��H�Mz�5��$G��e���y���W'J����;:�}4�C�LC�P^f�6�� ��\8h����6h�����g�&��(�������o�`�!m�x��2x�./�ڂ�R��8$�܄"w�8l�#Op��������H�R�e�+�����4��F�S,?*�ʠz&\�4�u���m]�@��euENK5ԢL 5�Ͻ�.CH�O.�WR�<�,�Q�H%*Il�ұ�U�� �7즖����P(�%���}�*�*)��o��O-�����	/q��+�u�Ǆ�yU���z�Z/pry\}��)G���/,;@�g悏�r�^^�D�"�JL9��w�Ӟk<i�7?�M[�%F #2�V�)t�UV/b�`��YBn)6�7��V��:��i`��]�Z:���`�ñ���؜h`ҙ��k(_m��c�;YX?���њ���c��#��s�&����qr�;�#^�4".S"��џ���_]w�EM��;?Jպ�Mj)��.�\�ŗd��'OS*X�a&4�$��%V��.�DR�sY�����{\łGb��Q>q`���<���Y栿�NZ��_TFH�#�Qo!b�\�{A������JHzB�G���%j��2@�����D��r3��q*����=dc×�C
����+����$r/4D���A�6y�_)���~&:x�JCa� |b��^+�i��˷Z&��l[�����=�a��m� $���

"���Ę췹��mږ7��`���m�{�9\�������:�O�`o��3��]��O乜�z�aT%PA˰oۥV��Zkoa���x��&�� �k
X�	��߻Fw\#$G݄�"��u8x�q��e�Ȟn*�SH���юp�N�4�yWE��9E@R2ك�! ��э�(�'V���0���0\	���ŨT�FH�
?Ǡ��;��^g���wZ�M@�uH�`�n�����`ا�/(
�[���W!�J��?�fX�W���+�7�>d�P`�h�N&|�4&t��hRD�E�����6��]��&K�f��Nm����/B�ϴí��}��`pr� �w���;/�y]lW�J�9����g�(�DRs,����s������Mdk�"�>��P�,
Y:S���G;1_�>�ސ�<�S��8�$�f8$G�jS%
n�!�^��Y���7D&+�����,�-��h�������O'�����Ft|�l��#�&_��C%+_%3,Q=φ�V�
�n
�!$�+�	������T�ݗ	��(�@\[q� 3��ԛ`�-�:@�x�~v�Ւ=ý�&�w�� �U�[��ࡴ�
���#�O�����~�L3�)�k�/��d��f�"�AnM���d_����I:��Z���~$�JQ�$�bZ.�̵�a�=\�&Y�5F�a����.0{Ym����#z�q��[������_F^$){4¼tc��ç����/��B�_A��eC�~�7�}�D���7L�x��ɚ��ʆ��'�i���ZL8n��z����Z���_���Saʸ�s5~����nC2DSgEA����� T@8�D�y��XC���s��G� #ЁdW��`�������e|ۀ���ulz�
K�}� ��pI5{5Wŕ�h�{`�a{ik�.�"�>�P���L�*� ��T���R��]dW�뻱N�S�P� �����(��nG�M//u�3������(��,��p�_�m���PoN�(����c@A�ݷ,X΋Xq�*�R"M�c�P�ђ�K6B�q�&�P�|^�;0Q_r��^�w����
������'o@a���H<z�l���$��O|�5���ߣ��B��D���OJ����:��G�bʽIn+����Wx:wZ�m?"I�Y�=�+Tg]�E�ʊ2��sJ�x.��y>dB�j:0�Į%�L�w?���:��-���?��:�SN�S��r��}C���&ž{B�L�)�($�`[��Ly���j^h�3�~Q��4����4�� Xu�iJ��{�X2�]M�Ҕt����(��-�{��hP�^h�:�i�%bX�,��Et1��G0��Lh;JKe��$Z�t�t����I�_S��'����o�c�b`�ow��<k��F��,�6݈�󫼅�Q�h<�Slt愬�_8���`se��얫.P�Ǻ/��%���9�|_��N��!p�gI��=Q�}:(��;����t��C!�4�Z�-�����ë��x�mC/���Z���3�]����c�S����~Ŏ1�~iAh��+���g��>I�Q������ z�W���r"���9JA�F�N�a�`��'��>�=!��
ֳ��P�ۇ6ʢQFtuE����U���Ly���c\a�Cw;���w��>�9T��(�ƽk�<VĐ�=����F] �A�]���.��qb!�NWұ�����F�jpL�/��(@�k(�ű���Ro�
_rB,"4��`�"�g�#:��
*�Mk�s��YFOfge�C�\�dg���j}���?T��Z.�f�� Q�E�0U�y%�#�7�OL����1�ԋM@�����m�2�11?c����?�M:��+��X*,�w:�AM7���X�	焣�^+�(����
M��+���T�gr	�E��-b�%��y}i��e��N]\�#$CW<t��n��4��i�P��ah��ty�.�sV�G
�	��tS���ɒ�1�r�ZF%�Rɶ�s�R�f�������%ru��@�0GC֡������\Bd��\�!���䢮N���WVSq5S�m����h�u4���UI�.ܮ�#c�תZ���'�3Ӭƌ�5Nh�ݡ�p%�5[����6�>o6�ԕ$�`�:7�nW�������f��s%��TC��Hp5x���U��q[N��]��8�F��ˆx������uO�.&�<%��6��q��F����#��*��ҝ�M�3�i�|C;ͩԼ��\�e��xp�����3�y<{k���!s���8��"�@����S�$���i�n3��r��H�9Z����ڕ5�ϳ	H|���"��{��Xg�87oI*;�b��sG��Fd�c�0Z�̝�������rk�����A��77隷F�$r�y��跕�k�jE�WM�Җ��Z^aA4��$*6�L�o=P��w�w�"%�6�>�q��m���MA�»����YcQ��@��Z����*��r�s����n�%g��q��!�5{�n/�9v����݄�$�]e���LU����<��Ki���,�������"�&�4� K�6k��`�x��`v>De 8OZ��gv�6�/����\;I~<b#����C�\l��g��]gp���ɝ��6�%�|�c?����zM�W�r4��L�X<PI�Ww�u<7u`I��hT5��ִw�~*;�lg��O�F�w `�~�����F��	�������aK4ȈH���WT.�C�ؐM�k7I��a��+~���U|%�V/��dj���-:� kC��[��u=���)�4���j�ח ���0�y���c�z��JEe��]�lEd"����O
&��[̉�h��0ZKjxw$��6�S�:�:�E:fK�W��y���]p��7��p�e��|�oΌ�硻7�k7�2]���?rʜ:b{NG�OD��Iv��?б�ax+4G� <���7ˀ���`�7���}Nsq'����a�uF2��=?��'���e�ˆ	éZ�]t���+�$��\�>f�Bف��a!-�I9�R��B~�z9c�L�:��ŉ�Ut��W/�����HS�D��W����OM#��d�S�� -)���l3�H5�>���	�,�<��9�ʾ���m҄W��%���`��D�������6!��j��
�&GE�� �kśc��m;�[�X"	|4_�|U�8B�޺����(�jMf�^,���&���1�{˖Uh�s�q���39K�d����Z�j�^~�'�a!\џ�ӵ�*�J1!�Z݀�xm1H�c�}c27(ٔVm4���>X�C�s@�)"�&��Ư��1,�S��F�����U��ߣ���)8�U:!ؚd��/}v�0$ir���J�®��yCc�廏{�l!�Rc����/r_l�P�M8[�VWdW��$��]��ҸO�S�ݝj�S�z� -l� �%H�阺�O4�����,����*�g�*�89c�M/"���@�q�� Oa\����0��>��<�G}&�jJ!s��D��l�GR��/�`�O�WV ���N'�F��A��
�����\���1�	aB�r�^�R��'�a3_SGc<Un��FˮV�F�o�������1zUڈ��s�k?(�(%x�{���'j#Tc>K�m��P(:�9�êdL��JCC�u����!¬�Vd�[K�P�pH� �U!:T9:x}�4{���IE�!�����W�n���Y
�1°<&)@@���©��C_����/�	�V{H��2b*�Hn�T7^�+��*�R�O��\�8&��Iq/[�p@�Ŏ������~�H�v��*�K�Ȩ��d�����b\L�Y}J�؈�����rQ?��Q35�`�MI,)\��ö@�F�^�������K�+&ɨk�gs�0],�m��+��AKT0�h�0E\�)6݅���H1Nd=E�����D<<Iɏ�K�$���%��Lb��<�L����{9�m
�t�v������8,�_�-���r=��Jx�{����~
zX�1j��L"H��-W��d�CsW����F0(Ńa0_����5��^�M�Y�c��Ӳu�+7XO��~׌�Q�DJ�G�ՠ�����%��ذ�$��I�"� X.�)[�I���3��Z�`s���R���c,�=�qZ���9a�{/gJ_u���|`�.��%�����얹6������ە8����0����!j�^Tf��ݠ�l���/�n���m���6:��8j�Y��C�)��D��j��>%Ʋ�B^�:��3�X�7��������tS�5�'��ε��-�
JlLoLe�҇�A ���@`E�o��c:W�{�%3��yܧ�g`���C�ݸ�۟�G���̋d��i��FF����[�@�:!\NNn��(���p"�b�qa�*Ք�|��Ԧ�L��Q��A��7���.�۲�H�Hc/X���yOy��y]a��F�X���l��D`L߿ur�1oGV�����G�l�q��L|�0���U>]q���]8�6�s�>�rd,�j�X>k����ܘ����o��?]��N,�E�R�0,�D#(��^�I�*h�%m���Uk����$EɃ?y�$Q"��$ �;:g��k��*V����CV�_����b3��Y����7�M���꾉�}��A��;�DKM��N��0�zo�� g�_:*ǧK?B��+q��������/���`���_�*�����҂�/lo訫Y���Jp5�ϝ�U��y;TkN��'��	���2Y�!�G�K	l8�8#��fa8g��+K�+�Y#��/7?�!�\�S�p4g;�^�0��5H�<���Ϩ��x���_tʛ��br�ϔ��,�^0��-'3��ҏR�q%{|�԰��D�2 ���1n�QĻ������]��6�9`�'A�M��5�{euJu�qȆҦ�������o(�:��:(O��ئ�V���eU,e�Y�t��./_|�n�����2��A��8��R�@ Th3�9�ᅷg{�i�z�n
�#fd�����@E���o��et?(B��P�x�R�?g�?^VT�����Q���f���]w�J�n�m4o��L����:���i�5���D���˝�{8=��^7�ϰ�2�x�4����M �E(�Z�O��
m���b�����<jJ����L��>F�i���<-�2	���;t�?�V%���`�KJ�R�������4E�������ͤ9ǟ��4��LF��ٍ x���5X�>��� 
/���h�R�fKp>a3;�6da��#��w&���cY:Ԅ����=�Y�$�[n�X��{N�\3Y6���EEr��l�j/�T7�M�$�S�4��lO!p�����#|3i>(J�"��̂�ʐ9���9��w�1���i���n�d��=̏�����Gެ?+4��׊���7�T�B�cX&`��C��o�W�d������+I���݆��J�S��X��t�TM�Q�}� +�Ȏ(ę0��#V��SvWfn}�4�KS����r�k���qY^ҕ����-����fP�N�u/-�
Jdb�.���	��p�u�*�8/��S�[�\#!��=R��vZ�OnA�]��
,$r$�z�UeJB´�t��"/�lp~\lc�4�����ݛ�w#i�Lg-��j���e��N|�o��Гi�t. ���|�o뾾nsı0��-���ףɄO)4��QU�b4��Pc\��9�����j���o�� o�+� ��U$!�Z�0P�S �=�w�%�m��]��Ψ�_�:/g��l�*�,�[�YO��?����L筤�q�a�&B_Nq�pE$�\��� �dS�5y��n���4~k���x�y���t����h}2.�f"7��Q��T �M��N E;φ�?n���5���;>J-�M�ր�]�3�)X���	���ӫ���9@�*4}"}��-��^)��L�Z��)�}߽}!8��0k�(+���0�����I�@�u�3��v�n�==s���
;�!�CV:��H��Җ���P�fwT@רy,�F�b8� �����R��m�-����.��0�4�ch����yA}���U�l�:�:���Q��4��=(O�6��}�]�,�E��)�l�G�zp�
y��Fm�BB��׈U�\Փ>4��D�9_8R�'��E�����6!�W���o�l�Ę����ťv��h�o/#���C\���K�%�} ����V����n��d%�H���������L��M7�䌬*T~O�4�J�_�[���4��g�ϊ�[^N'v�mG�
�#� ��N���}���u6@����Q+9��l�ϯj�V'e}DB�1��+��Q�\���!���P�i�~X#S-�*�)�#��0uD�	/�dB����v�I^�m@�N�a;X���Odz���)^S�\�t�z+���V��b�P=�%&���@g�f�_��Z\��!c1�JۿӸ��!���~�?h ��HM���W��pL��S.仜�Ad��#f�f�C?a^�n�d%Grm����% ��8T����2���+���{�������44P?����>��.}���n��� g`�]��_��Y$���N@W�M�������]���G�a�"&��3�I�,C7��^弍��������Oy=sߌ@�n�
Q�>��RC�M��:Ոꬔ%\�@Z-�A�P�~r��E.r���,*�)�Ȱ�r��/�P倊s��{��0�ȗ$1���}�C ��T�f���&��+ɿ&[�Y�G[Q�4
f���A�4b&Ɨ�3Lnp����=���,�b�"�üims��g6�M#���] bބ���j~)�dD�_r��Ѯ�Ql���l>�e�?��[����k��롔��"��J\�� ��l	LWð1�Ub�!K�\X�>�*�p��%0�j�3�t����<b�W��9�~β��s>o��q; `�_z�97�t��?��|ݾE�kiPO/TF8��0�d�*�zU�$ngi�)��X�Gt�%�?�*��j��7Z{��B�*bCO�9f�И�f�@@aB1K��u����!Q�3w��om�N��w}t��Wߓ�i�Gv���X|y�߳HG`�۾��fȉ?��Y��ѐJ�wL(6U�˸[��	�#z�+4��
 ^ϮŨ�RX=Y-�$��7ܰ�x;2(�4"2��&�⒘����6�����݇�EX���Њf��o�*��<�DVi�|��H]�����G��뙶�
k��1.��J�������iY�<�J:-���;4'�/1�#' 4}s�+zM�I	��MѾ̪>���`����/��l�C �6�Vq�I��Z����`��k��j���u&U-�����ꩧ�Ut>Q��1J����y���W���9	�¯Z%�j8~�j<:6K�V��0¸፩�6��B����s�
���\�M���b�{�����C�8�F��O���;jK0�P,d��S�p�i�-��4�I/'�ķH�7Y` ��,�`_�1�W�r ��	�x	~
��B����!D��!1�C��qu;�����O�F���}�K_��V� ��k��͠�'�ח�6Cۊl¼0J��[��L�j�LE��x�4F�9=P�y��N;���K?�C�<R�7�l@u�)����v�6��$�8��\��*�+Dh��7q�D�JRte�Ġ��[�j�^7�a����$y
��I�:Ef)/��^�.�EJ@�c��@������z�������	�\�(]���#�wkr�ͣ�U9L����%>���d7�2Ù������TK(����(;��p|6�P�7ܵջz�>�v����[S�����#n@�y���#�����`E8�׷}Z/cM�k�+�����R�w��Oh��GB����VP`�����3��3�T;Ö��{v�	������0�G
C��H,�g�'ض h��Sh��q��0�ԣ�s��xv�e�j�'t��o�^"����H���P����Nz�~�K�s������=��vl���'
���U7�)o^ֆ��xD����擉ehj���|@l��KlzK5�H0:rƑd)�-�ɸ�F���u���M���~�Y�20K�����Xr��*�8�H�>XA k]����F㖕\ne�p!򳌋�=��6,����]�[9t�?���"��ΜK�y�զyt
�yjuì��^�6p��-���ly�_]�7sIS'Z8�m�v��}�������X����+|�Cj� �/�L1K������E�ш ��j�݈M��JP�>�8�s^���nw%�D�:M�����Ƚ�Jj����yx�j�	ߪ�h4daVޫ���Ca{'U�Ž������6;�C��=�WN>����7�ic�o�</��{�����})�E wt^ӻ�8{�۝���-i�h��lڧ�|�i�8��E�B��ݱ�6.���VV���l�q3��еB���U�ı���8� �:~vV��z����Q���WG)ia�G���vbE~ݼ��G=�	Z�N�)���ǰٓ�RJh�MG�'���W�Q����ܿN�lƧ�����H��T�O�F<v	�'���K?g��/B�^,]�>qD֗"X>�L�g�C���v,�ݩd:�à������r@������Vu�Q��x?m=@@�w�s�@��ܦ_��ĆG�/NY��M��D�S&ʉ�M7���5��w��{����o���m���*����{�������<��V�Q�*i���'8Z:���a�?gf���E���U�ٵI���QѸ�]Ң�����?�(��Ր_�ڂ8!^Lk*Iր��O}�7M�w�8���� ��/1=�)�ז�d�Q����Q��qC���4ّ1?!��oF6�p+������S�1����n)4R�:�h;%ad�v�vO�@�(�b����A�i�d� N�,���OM��(������FD2��U�Eǘ���Nz�&)cZr���Ǝʅ�s%�w*�6�}P�w~Nk��AJ��MGj�i&G�|�Ņp"(�lb��;�V��K%v�cI��N�t��͢R[�Ď/�/��Ѓ1���q��⷏^��̥�my>)��֐���G��<�R��މ�\ޝn^x��h��� |�z��E�U����<��m9�\}�z3O/o�]pߴ될�������R~�ݠ-���g>#��s����:���Epnb��!+��^k�Op��2d�@$�'���Ś�-�ԧ�x�&Z�qӒ�o~�A#����\w[M����D��YDc�m'\��,\�}v�a)��N�G�W4ap@�P��T[�7?tM�g��9�x:�g� Ɲ�����&���þ�]���I#
г����ى��3���}�m"�'bˊ�!>��՜IMau���G�!�h��PD_�ݨ&�p9`H�rͮ��f�{s�S(:{�e�K1G̩�kf�]`��A���1;O�1;��?��r�^<��cP���7�q�ҋ��F�B~�:W�*�
>���.�Z&���"p�/'YXi�8�t�u��5�A�N2�Z�	(r��� 踟N��ъ�q�)��/&]��ZaOB�J1�c��s{r�`>9]�2.h�BH��=��1��u�H��%�^�j�e��%�O��i����_�:��`Z���Ɩe��X5�v��0G�؂��1��8����b�9�پl2��F��8}gEƴR�8��K��v���s- b>\�  8\<�M�*t{���~@�m	X43�ڄ��~���H�w����f�U
:�k{8�Nf�7��ȋ�={YujIX��h��1�oc�f�_ص> ��0�.���,���a1�{q��N�%!���ig�|�(g�0\N=W:�dwdw�s�Yw�*��q�&���zc�$^�'�QN����)����ۧ��~*%F�eH-�	��U�(��k��A)�m�V(��8�o��D_0oJ�z#9).�*�+�re\8$oe�߳�����}�>��� 壒�H73���O��WM�daDӄ����)�I��Ղ��������^Ihԧ7F�P������33�Y��,�7]O���E@����?��tp���{S���-�o^�ۥ�����te���%�o�b6�/���*�{�L'K�S���S	'/-�c���7L����Dq�.Sg�H�����N3�X��>a�b��gk!!�f�l�x<Y��'�<#A�Q&�v-��=���;u���f�_��\u���8�������m@��=m@VQ8�D4,�)���Ŏ�U��?[�}�٧'I��������p+���o�D����w`k#�����iE� ���?H�'�Y�4�J����+�W��c�Z�����3�V��y�wE
Cة��޳����'I~c�
�M��U�J���w�j��M^��QT6_��>��,pJS��,����vGbsP(B_�T�h/�{��d��g���w8��^��W=d֗��4x���O��ɂ�4(���2|�ۊ��kA�I�W�	"��;k�KM�/��G��l"g���ߧL>$��l�b6��Á'D��5	P�TW?v9�����@? �~��~H3'R`u�=�b4j^� ��-��E�A������߃&����d �v�������n�_Կ[��G��>���w�֪�q���3>%����7+V>��i���Ɏ����yy��E��L��![�,�Z
z'j\QD�����H6]k��C�>;p��M����ύB�Kg�!���I��ҭ�aՉ�VR*�N.I�֞�^\,�DNV�7�1���BWC��C6� 7��X�%�O�(-s�@Ft����]B�kH����G��6�/ґ�#y��� k��P����ǆ�A0��k�>�Y���$b���y��[�}���߄��ٓ�`.��������ڴ��u��8�u%��}��� ^H�T@����Q��9|�>/���QL���ΐ�gܮy��;�Q$UǨ]x�f0�aeU7���`�#r=�P#�ߦ��'�3�����a(�X�BW
.�s���N�4�U��b �W��RC���/����l߳����!�y�|Mv-g1�2��	7|�٭�]�5W�j��G�K�m��B2#\vO�r����W;Ţt���F���b*��.�婰�+�؁Z��T��׿��={Pn�f�F��I���P�����q<qp_��p@��:�#(贅Fp+�q5�v��JW��oC�˥Fo~*�B�������/��Bp��	=*'>���>�~�{ñ��4�����ǽ�?-��R���Z��s�$���
�|%#[��%wh��J8d�b#8��-� ���4�d��K�å�W`�cH�ǜ�隒�H�F�/'�p�����9��������#�z��f�v��ߝ�ZB�)3�S�ʋ��%=U	�A c� h�`�^�%J����U��G�&E
��k��:��>l��O4o�2=)u���ͥ����+��}���`w��G� �:�H$�J �.�e?jR]X�|�8:Y("��bd�uQ�]n�k�Ze���n���{Kr L�,�aӬ�����Z�Q�x���Y_��\������9V��F/�\mQ�Z��N�I�n�n�*%z �� /.��I�:u�%�7W��D���=��-S�<{�ؑ�UU7{�R]��A�G����C�N�$<�j�@t��2�k�9�;�ޤ���؜/��+q{	��N@gx�+zLE��pJ�Y�����*�`1�-<���h��/�u�&�&�gR�*�;R�N����HK�'x�� ��O���:�zH?�iJ��i���K"�m�h$���K,P���"�N1�R@��.i�J{t�7ڏz�^|FU+�1��G�K����� UL�~�1Qtbm0J��,�P�{2��~�tV�[>%��W��\�:���UQ�3�H��z��A()�j���I�������s��P��aO�N���z����ҭ��n�$E�Մ��n(;NB���N�K��7X���㠭�Y���l�ww^��s�9ԯeU x1!�}���R:��{ƪ�}��:��M!um��ˏ-0���"y���l�W^��P�9|�$��'Ma[9G��e�<�V�b*	oJ�N����L�e�m�̀S�]#6@�U?�3�8qG>P\/�*{���"�1��l�abꋂ��/�G��n���57�
�WWy�ى ���������[Kj]�yD�i����(��5ڭ�f��wu�y�k�������n��8��vY� &	���!��l� �#T�+�i���r��z�<wl�E_*��<8�&b�G �sF7�Q�����X	No�{��#�5����&�Zun���V�W�~#|��?�̫�M41.�J�[�DF�H{Y9���x�s4;S��AŌ��`W9$���7bYC�2Xp����]�������OZt5��~٨�}Ex�
��)�	�O�0�/ʋ�b�G�|��o�E���?�XO�'~�Y�g@#�>��p@>����iu�;�*��?�����n�jR@�ϔ�{�	����/�]�Q��T嚈�Az&v��ڋs��� ��Gc���6)n�����:_�D%�ۇ��>�B���`d��G=�g�m&u��x"�A��C0[ �8(���ڹ��7����4����nk ���Y�،3����;�r�Ά��]�i��<�-�t:C	�(ڄ}3�I�}����cx�ύN�p�;�/O�[%J)���J�oF�J�ݷ׊��� �8��k�fn��'VyD���"�j-��`���(����_���=��ID�=��Y�����Z�08leR1�����Z�oZ��ĝpc�UƏ6�����͵r� �/�I�����p�-H�6��60���|a�:��[隷�~M�/~�-P56�-4<k�_�֤y(ּ�.��X;�6����Ub_&�Ɵ�����d�(%�j�k���k#�R��������qlRg�U�\x�2��huN���?R6����C��Ǳ�(!2�R��Y�S*�G�RQ��c�A}l0�9׽3�K|f�:!�}4{���Dk�H�s�] C�ͱ���'��@b�����;דD��DuV��X��p&,M!4�u�W�q���D��h�};�׶L �m�~�~Py�<���c!��݇�9Һ'�+%�%��g{�T���#��0�����%���@l��l�����&βo�0�M8NN�o����G2	z�蝎҃�E���j羅����n;f=�(Ke �j]�Vv?�.��,���CuVcĦ����z�
��1�᪯Ȗ�$��-u3n$XlsH��]�L*�h~�=�ד���> ����=�Le�e���OqF�Qh�&Ty)���d{���;(�E��D�Q�Pإ��h��i���sU'�40�?��.:v H���:�s�qӡu�8����U�uK�9���#VLm�Ҙ ie��d����#���=����9�HƲ҂Ȋ(�� �#����r�~���a쨹4��&J�7Q������Z�Z��t��-�:>аi�9T��];�8�D����e����U6yr�bX��پ�
�D������5A�yL��@�]�^���Ɍ5�>d1~�1[��M����?�~%Uܙ�T{�9��!�fd��-g�}�k�s��zg�l�X��"4�J�t5c��.���,��t�yS m��A��,rwVi���.�`g{ް���ډ6m��Tٍq�i��
^E�N�{��g����W�����
BkŎ��"��.JUʜ-���3H�:��~'H�i���k�7��;+����m��닋�r@}�v�#<��|WW��j�V.!�n�o@^��}B.�:ն���$����f�I;�Hj,Eg,4�4�������z�G���FM��+tP��m�/�k3�ģsj�B��_T
֏>N�À�|r��^��m��e��^m`���~;Nա6��N����s�E/�^��Q'�*�'�!N�BR�J��h�>ᬅ�(��(s�~�h�+Z�`ޓ�aj��^S���?�}�/��Nn���P��h;�ԛG��3ЁM��r��H�x3\j���]c�X����CA<�[#!��q��@�p_�)���F����!7@9��Z�D�n�=j��h�ϳ��W�UZ�#��mZ�J���� ��&�Gg��g����.�JCrW�T���>��X�����*h�U�3����{"���XtU�B�� ��p,�h��!ǽ�(�
��Ԩt�4r|����֛{B����O�Rx�q���5�����s^u��]�7�Ph�1 �NOS�8�x+%;0�䆥�բ"���JZ#�3k	������Q��6�|������'����Ɩ[�,UF���Q�*N|�ό�$g��(�9���ʭ6�Fc��p�_���NM���NXԐ� �'�9�cH-7�Ss;B�\!vG��
�P�����&n%6rڵq��Ý��2jy"�d�P[a\	�=�}��`"���U��M�ID�cE��l+�� LxQ)0�G"��!�5Z�%�*=Q�pk$ᔱj�)���}f���W5s�jܦ	䮎t
�nԍ~�A��[En�>��>>Yu�Y������p��n��E.Ҧqz̴�j����!���Tdo�)k�J+�<��v���t�HR�T�]�����y�J?<2Ƨ2���N��r�+�"�c��A��m����?�S�l�S���Pc^���O�ǯ��w��OJ�T;- ����u���T�	�o��ʜ�]$<�S��4B�R!��=�h}�I�-��o����35a�-ͼ�hS�8����EO "�W��u�lf:G����^���"X��bW[�v6�z��;�R��;�4��#�^�T��:�X%�j�V?eʵ��aR�/��)*�O�3�ci�q1c�}�bl��G��U��{�д�w��Ɨ��.���5��[�Z��p���eg��n�''���Z�	�S])�?��h%�p�3���\�}g�;ͭ����b����~�����\��Qp�u�6ﶦ��E�ƥ��U�~�0$f~��HMs�]�K-e-�QB�u�P�ec���bmY^'p"�
6,��� Ks�/շ�P�����Յ�������`��.����Y�c�a4,��l)��
M�@���)�P>T����	�BG���Dk9%�O�fB�k�Q\�� 6�9\��t�5cO݋!�>�f�^���x�S0�u���݇��n���g�7�"1Q�Ӡ���k��ryTDp#��pt�wA&�I�7���6���x�K��Q�W0?AQFLi2.7�2��
J�&r6�\��CPP��y���U��RY���b�`��XB\Hko����:1�"��%�g����/�햦X�Ҧ��'E` D�_�� �a��%Ą��w�8��%�d���O��7�5�\Ҙܘ��9�+�b��WX:�����\�̩<��	mǓp�#(h��E{-���2�D��4󦺴�>��=�1J�����v��Cg�iE%�LK�J˄&��c*Ty����N�=ZR�N����M�7	�Zも+ו�ϵg�9�F ���T.����s����x�	3�Jeޜ�Vƍc�R��>[o��킖^8|�i�vh���wYN�dMI���3��2,�+]��<�0A�N�j�oj��u���)Ȕ�WN�}V�b�-��Ձ��u�hm �����4�!�^v�������?x<᳾�K+,n1 7`����O�.V=g����ˬٯ��9\�=�}�GC��d�G�I�$�g�@/��V\��y�u �rM��|�1o=
�����ܧ��f���n�y����k��(D �4k��W�G0�Q��� 2��)O��=���mu��H4�5���T�������z�r�J$.K)�C+�a���jJ=Ό�����n�:eI�:�9! Fڧ�\>A�?��eO��Ȩ'��į�+F� �E8�ԧ��Vp��B�n�~���X2��v�s\ ���Iȩ�]�q��.�����@yp!��#A����0]��'�sf&S-�3�8���g��)i,9�>���]�`����N9�C�kڷ_ctu��x��U��.ة��[�$�M3�B>Y� :�����26O �;��,����nO*m�����b���}�1�P���bC�s����Y0���qO�y�몮s#���:�����A��W�R���U����<���q����EMlԘ��n�Y��tS-���[A�]��n�S��c���p��w�9�g��&�+�F��)�U'��J�@��q᧐�ᘳk����b2\�"��˽/��G�;:y\caK�`Zq����re��/�1)��?��Ko�����ݝo��o�e���`Yvq���V��	�0�n*Ӕk����b���x���E[��J " ��7��/�J��U'a]0E���n�����#nH�yz�^
�\�j�F5� !r9��Jz1b��1��GG�û=}}���C��l3�Gq�/5�"��MĎ�
�*���?Y�C��|��Zĉ�,�A����̻���v��/���y;�Hԛ��+�P�V�[�%��id��0��qjơ�z_M�j�V�z��4��0�^�P0Zt�.v��fx�C�C�:�A�Y�:@$g�T&E�,�(���phA��<
��Ź���00d�ċ�Ɛ��~�OOL��qR�6�@����rQ:c�N�}�I?�-䙕\�T���9qX�����y��m���&����l����=~�o[H]��[ݦ�������k)Ըŷy���4̙v�mo�9w������r�I�+��<�~C�Qu`��nX�a.�dWX؆���T��eb} �4�1�)�����.g��Ȕ���GDr,,��Մ[���Dhb3���0�T���ne��OyO�d�b>é�͕��2�������Q�!W�{�fu �5[���!$��01��4��%��_IN�%}�d2x���c��h6ɣ��+��t����g~�1�<�աN3����ᲁY��qeL�^t:��Ja���*����z�U��k�qt��V{卟/�	bE�wL{)����������tm} .��`&ѝ�������e��JU�p�1=6��Ȱ�Kf�:�b�݅Xur�Ȥ�
>���+�t��S��bW|j�"�^�m�`�ԹH[
�x>Z�N9���+��oM_T~���E�n����\-�Zm�jm�Vҥb�koM�]�ǁL*�4���E���.��Z�2T�oQ�� ��놉�+��Ό�^�}"�
���:����Ԣc���Ԕ�^��a4���Nۼy![^)ZL��	E4Pe!c�*y_�Mг�G88ŗ��%H�6�E�� n���m~�$�r,wWɾ�>V���e�m��U��G	N�X�`]P��8Bt�_������q�K/����4m'���x������τ�^�� vn3v6q�2�B+�"�ԟ�o�� �ˆa6̏$�./��L���[TIdO'�fC������T}.~�N�U"3�Ǔh{�Q@BaiǫޘW��_��s)iE���7��d��k�h��]D�7����C�K7ʻ�=�1��\U=�!�=vLb���$3q�L�_��5,��+�搦g ��HB�,�8m6#���,�a��/���L�y�/C�d����A��)W \+�c�����<ɼ�v;���K8n�fJ~�~���-�wp��_;�\��lq&��L�[�#��Af�x��~�����*GU�U�\3R��x��e�`��M2^H��Ѳ�Th��B^�<���w�R�������X[	m��Q�wA����(�Krt��A)��3JCޤD=�����p(����� z)�J��"d!�Őtԁ�\qگ�6�G��I����95���\��Sv�~�(��ʨ��V�o����������?SQ(/���)���d��a(]��퐃��*�3ʳƬ�=�y�����;Z�hD�_d$R@�y�����tR�.N�Q�v]�,��\��b�пa�C�6�wp��'Ɩrs!Ci����\5��YS��B��q ~�E٨�V:L�)L��d�Ǖᏼ/w�T��)�SS�h��{Oܿ.t�!~����s}��k��?��ȭ��f��X��< ��r7��߃�6H��+ދ�S�ᵡ�DJ��ˁI�9�¤{�A9��t�r��kg�,������d��b�:�ì3;�� ��3*o|���,�c}�噭���ÿz��:w7A?n��k��{u�m����"E����sO�UĖ��c�Z�TW�[��iD���z�̌h�G;�D� �o_H� 8� �E�� \�V����|�BYEee��t�v�yBw�T�3��D��:T�d.�sG�?1�X����Q�h�B������)t�'���(F��if HA�w��v�	x�3~���}b�&�
=F��cUשt3����S�ԃo�,K�]���=V��D@���eP��
��v}��k퐊����;/�q��onDt�#R�1?�wB���U�w cH�kv�+����X:���3�Ҫ�p�n�����cҋ4�2�p���IۭE��Xt�>�`��n�j����!��۷�}~#_�9��BC;p�?��ϡ��L�!���:¹��&t�P�s[[���u�x=�Y�R��18H�3D)���cQ�k-�z��E��"E�_����Q��hÀ��ׄ��{;��O�z� s���2�9]�_C�ϥ$��.Se����wu6��rVS�#�h�@�k͵�}�)���|�m/������5!��`��9���zb� c��/�����?@[tI;>s�M��E��S�5���<�+��6�O����@���9[��E�14�
���Ť���ū���*��%9]
��zT���5�i��5���[|~C������"�px�=N��eW�@�q��ѕ�'���Ls�*H�MbwE�~r˧���w��^���(�u�o������+�R�[UڪM���M&�W����ee.��Y��F����fc�8R�&G�� �"��!PkF3~YJ�8\1�Z��ݴ�x����&��oj
�%!0
9tM^*	�M�:��;Y�k�N��9}v�|�D�#m)e�+E:���F�{�ł}�����7N��P�MhH��:��3�����"QJ���ڭ^@��mu�p��8N�Km�%G6>ü��k�_-<ZD���u�g��\����W��s;R�z-���X����0�p�A3��".�]y��������GlZ�����O��PU�M�	��v��*��e\�^���N�ZH�J�X8q]�SvE�y�r���!��%]&G��2��1>���M�����������'��KKDb�UP��Ճ,a$'�U�f�TB������[S�Xq-�vOe!A��G1�F6A�F�Qb� �y�7�����Poˈ�rx���ܓ�-��g4�������+9�)���
s�֗ׯ�����2����"�t�M����;����y� U{E�4gM�r("<sy��Ϥ�%L��3����A��'�?��/n�R�'o�Ŝ1Q��ŋ{d/_��H���R"��H/�I�_�<��
>��Xk�������#`k�R��)Rk7�ҋge-h6H���`�ߦ���6`�Q򞥅�f�j_�_e���1�\�ŉ����1O�0�R���תS�BN��(�ǰ�h"l����+IqK��W��0 .����z�sa:�f��ba�P蠥�L�z=k�~�c�\iu�$w)�`Fz�7����>�Ɩ ���5��iF/�����*h�ԩ��=_��5N��x>p}L
>�p��w�k̐$+�	�YJnj�eCU_�T����L�Q��Q�AN�v�5~��؇��O�=���3��n���K�9�7;�61U$ƴ\�
�n�°pL��A1B	�)r%VIm�3��v��}��8w߈.��a��նҙV-Ò�L�����y�@"�{.�ŭ����d�j�Q��Ovއs�h�J�X�C���)k���r�4r���r/�:��,�ЊkK�2y���i�JG�`Ĥ�9A�T�G��HӋw���F��HQ��Jwz!��/� &�N�71��mC9Ce&Y�fF9)������I��9'�Q�;Q�؀ÚAfU�1p��^��>�Xu�
`7n#�Ȳ_,�Pb��@����7NE�p��Ղ�u����c�B��S�7�B��f�m:E�PxR�=����{��(z`G��;+$��z�7����-�Ĩ�p ���#{3�� ���Z ) ��ɠ��>�m���T%�m�~eA��yU�%8{�wJ����a�
w���ꢙ��SUn��/9>����B {���R] �++�)���ܗi����5j�/�w/�����:Β��5�"C��C���Ӎ��%h�� �-:�8���/�6�HљA\�q\���O����W��r,�*��%V�^g$�����u9��!ǚ��k��d!{��ˢ6)����'5zB�3�)=�<��]�@���`���o3���0���7���֞����}�q�3i����=�-�KO�o<��#���+M,����6mw�
�׻�e��|���[��䇿��-��}]έ���aw]�z��Ü���K��d/�.U�VZ]������FF_c<>��M��n����0������a&�Qt}��?l�A�&h�v���m����U�2�������s������M=Zfo�no��$~	�C�3$6�w�+2�Om
�|�\'���G68��P�j�-=|K8��$- 2�90h�z��v]�,>��V���)�����E��	dF����[6�+�n}(�wB�N�N��g��Y�ntm�ʥ{O@g�Rk�CL�@�DkLު�И�G�[��)6�p�ݛ�FsM��,�N�Ң�<�f�V>Ř���f������N�2����1�=�T��N�#ߧпM��vd�&���~� �*߯�b�>:M�Zs��23�I?ᵨ]��EWEu�wd��+ֳ�Jߑ��{`e�f��S=]0M��O�9���Ő0�sMn�N�x���J�B�F;�1F+�kGY��ĺ�T��?��� �RƘm��¾Ypڮ��U"�+q1wN�LM�fq(�|b�W��KL&�W =1,�D���>�yo-���<��w?��Ԯ]�Ҋ�B�S^_z���]�H������'z�%�����T����);l'�׌��	�9g�`���
���=#���������k���6Nm;�������X���%c�<3�y6�Q^��"^oٟ�ֆG�{�z�'�XF��2���/^�����]�O�Ґ��Ɓ��)�+�$B���8&P{��J�p h4�&�C���)�t�:�%�_��JG�~���ze������W.[�ҺN �Q�E�/��$�/!cA�6p��H<rމE`���sZ��n�h���o�JK�9�p�
�

�0�j��QT����Z��v��'�x��H��������elH���Rp�d�"l��[�|��W� ����g]�CҪ�pX�wf�5F�(���7�TAF{��z�F�Atg��<�V�$���{�/g���GIvyZhB�60��}o�/�d��w//��A���qR�KҴ�<$x�լ�T�cj��ۢK�^z�"cL*�v?�.'�v��M�� (=@l��c�0���~��,�K��n���9�*���� ׆�2���<�2aZl)�A���a�1��˳|�-ҪrUk���O4\�4������= 0\գ�(��ʉ�q\i��a�j����r�}���~����s^U2����p�m	��op�H�^��{S7��c���c�d�="b�9���3.��0��2Fr��Z�r��5�V&�sF(;�p۲,n����]��� � �r��l��|��}&��?좿��BJ"�}1YB|�=ۀw��V,v�吥�� �2FCOfM�?:Qh	�r�x]��`�E2"�����*|xw�X��]��!������e��V��N���T�|q^��-ڒ��N+ھC��]�@�^�%l=t�X����e8<���JRbbU��y@��M�3�9���)�J3:�c�csڞ��9�n�H�Be�fe]}��1�H/O��ٵ��p�F(��X ˣѢ�F�7u]�T}-��u�ɪ^{� ��س�{Sp1��=U���%�A�Ԑ"w�C���D#���Bo`h��P�8�R��bU�P��kt]y����%����t�Бs]�sm�b(��I��v�<;��RB)�����b�s��F�'1/�&!	�>)��	����K
��v|���r`ݸ^,�j���HJZ�j�l���t��%���5_w���v���^��I����k��O�֦6�L�4���Lc|�w���٨�`.��$��i80�;�Hbؠ�Z����ư#>���$�fu��M���K�u���qx��ǿ�1���V>��Nخ�`�%z8a�"��٫��F��{H��ׯ�V>/#�^s�*�3Vڀ"�{C
����(��YB�=!�Z_� ���=������u6^�-"��Oo6� �w�f���_���O�N��Oá���X�* ��?���¯��B@{�V��OGD���(���M��cy�?IOAFB'�j��K�5��
�5Y\�?W��$@ל�%�҂���obٵq|�m��۹N^O�<o��t��4l�L����Բ�m�
�!��p�N8<&�f��X�S{Z��V�ϒe���;��0S�O2^���Aa�QW\ㅔ�����%n{2�H{� N���{�-��՞&�lr�:���r	�<�R��.r�^���'��4�?�#P�v�V�z��,����9����Krt�ݪ��i��A�wʅ�f���@K�x
�'�~�g��G�oБ�^%``X����Xi�����b���o�=i����^����eY�:<��������d�֮�$]�o<"ϋ�͈��^M�C�����t�BF7�����4Q��[�'E^P	O����P�@�������ߝ����&D#(-t��r��f����p'啊���̅�.�y�S��~I����[�,7I���l�?nn��Q��oC�A�c&���Z��ϬDZ�[�*}��PE���eC�>W���V�a�������hsH�dR��H���0��w��S
�t�B�j�l�y��_Y�<2K����M���Z�ěO	7Б�:d������}B��J�f�֕?�@�#D�
�����|p�S�)��c�:�v�O�v�Z�NI��D�(�lSE��ۤ.�)�"ÝB��/��8��HMp�^^��T��G�B��I�:��LK)�S"(�q�LDZ?�a�0+����q���e��㢬�?���V4��@���c�V�q�hp]��j"h�zZXF���C�@�}~�z�����)0�)by�8쯝�|t�`]��L�ˏ�\c���H�݂Wʜ.$�7|м�1T��� g�~��`d��"̙|׵q���â�ՄT��.���1�G��^�Ǚ{�0t6�����&���@�Zϫ����Ux("�!#|�U`B!���g��Nx$��aǻp�I�q��z�T�F�e���{�ʧV�}�A�F\�=T����{i�aTLƍ�ن:?l��KS�w^��0w7����Q�����8��;ŭ���\�{�ء7mA��-�ڶ?��e35����Z-�Nw��jI��V�K,�~+-�P��M�b�k��x�e�\G�峐��ϓ_���2��ܴ`��+aV�$6AW8�&�/4�Y�<he1;U������w��2py�>ʼR�M��"b�5�|s=�k�_OTw<�P	�hk����a`B���<�\�۪M�T../e�\��C?��ʾ�㘑�C���L�����|9��`4�����S�Sd�����E�K��7��2�S]sĹQn��\7�]J��=���h!f���̤c!H�n"���?֓T�b���� x1{��`�����ۂs@JpC�-�#\�'�rS��Z_�~��]쑧Ǻ%����ǖ�e�᪦����I�8�-�F|��Y�i���P�v��2U�����(��?;���碤
Lԅ\���.R�{� ��Xڳ�/ۙ�����2��;�k�����U�x2>݋����d�H0B��4��y�����o��W8�������O2�7��1�����^M�(	��M��4��}�<c���;ϸ5e�e�rQ5 Iv��bH�h�ۂ��Wr�ͫ�j� �f�5�T��n���� ���\E��Bu~�TÓ�\cO:�3�P�ml�i픹|�ɬ^�>xL���m�K1���i�Z?�V!���˘��?������3�À��-��+ѫ�W���^o��������(�1��%�4G�mm�^K�d�����z���}yp�*�<N�aX`���H����xPW�>�ɣ��j3p?��]�����hAh5��\�G��(����^���qL��Jb�^ځ�j���K�Nf�G�AW������^ٴ�a��օ��`�`=D�O�|�lHJ���c���H�0`�J����.���ğһm3�+�� �w�4*(=��F����z%x���^��ГWm	^)S���WF�PsZ���U���hx��Ϗ�N�-Pl�(�\��U�K�Y����9��|�V�Ĺ��<U��瑳E���V�A	���Dp���^�(�=��}6�������Ӽ�tTe
������.�u���b��\#��{V�-�r
���%}+�PF�ևM�l���Cj ����8��zrQԎJ7P�T��M~�s�t� -�sybj ����z�5>D�(�v�u�����/jl����DM���q-�~����JwoEӮ[���#S�<�R��j�_׮��?����؞�K�����u�8Dٻ5�����9��"�O�����H`H�˿Ö���c��9��i�u��D���	`J�t��!'�T^�3�Hi�Աw���*@a�T��J�I�\�
'	Πh��%JN��hzﾗb�V=5)�{Y�q��`�Q]6���s�����#��=j��/�69���5L��쭷m�Z2�t7z/�� ��qT	��q0�v���i�$7����8L�z3sB� p����^nĻ.�_���[9�!Qhm��P1"�F4�4=���m�#��iCx���N��Iua�l�_s�d8	JJ���)����^V;���ro7�e�3��v����%L,]��;}�[�0�@� LG��ꋎ�c�3ɐ/nL來�:�����+���G��_�܊�$�>���0e�L���݋˟R��9x�H:�����@������I�ܗGR�\���)��@�cX�;n|Z5�E�a����\<x��9��zﾸ����76������2�swW�9�'A���W����g�h��8��3+��\B��0\����Ѥ�+eo
�š��eO��Y�*��^�n���PN��U90�x��B�4ς;���$˕��*��X�4�`��L�:٬t�/>c�%��S0<錸ڛg���d�};�ֲe�F���̓6����.�9O��Gf�H��^��?Vs�����bp����LѲ� �^��4��I\}�lX<S&��bC9�ݏ0�z��N	�y>Ǡw��ː�㡰�㽮Q���@(�ī�E[�b�U���Ho��p/���@>c�"������|Hu���;��*�_�9N����~fq�	�ӆu��4��l���5/���[)@o/d>BF��V�N^�`� ��?J�r)����b�ߙ0���V�V#&x�퉵��V�19I�)��-SB�ѕ]�?�#Ex��vj��~��byͿ�k]X�����"@4����^���ހ��%5�<��]��n@S��@�\���9UE.E~�߿g��]��ϛ�;���_�#�����zL3��7�:LG�K�NӁ�&�?A�7�IdY�(�Ҏ}�%G�=B���h����U%��9ać89�%�	8�~o
���F��'�0e�'+9�?b��k#��|�����V�XIh�P�r�42um�=[3PH�GOa�f���3�W�$�����@f��h���Cz���ЖH�
AV�s�θ����{k�y?��H�O�,V���]4�������Y�ŭE�z�"�Vd�_�S<�������`��/M��
"�輠F�����9���b����B1�ㅷ�A�Q35�F���7Xԇ���.�J���}-��`|Y+9�5y҃g��U"��ZH��ȑ+���
{{�k� %��"�Q�(q}BM~{
��jO/]/��^�Bz�Z���@���0Tg������d�GI2�s����=��Z#��Ͷ��C�;1I&��3cc*��G݀ٮc@h��V����B(���%n]��~*п'sw�`�ܔ"��� ��(E����P �Y_v���H��$�K�5�Ol���#�Q��~8Fݕ&����2`�<���7�x��?�9ծq����q�3y2
�ۀBf�z� �|���N�s#=r,>�AUã+5�H�6��YFj�V�]�s7^��;)c;��JpF "�H��!���6N���wԓSP=2Jt�\ܜ{���4.�jK����]�Fvl}H~�THkA:�h?Xi�pt�"���I9\�@Z�� �ܩ�_��C�� Z�t!���m��Z"[9�2N^��θ98��ѝ\]���A�%���6q�?i�AgG .0 
Cm�{�?��o���s���8��1�z&��s�u�m�ơ?J����d��n�}e�|��̓�ʣ��yH�|܏?���$!���-u��ɹf��1e�5<�94f��;��,�Z��c�>�L�����QUMX�6Z�y+'�T�ϗ��3-��Un`������OQ�YQ��0��l0��L<CF-��u�Mb���ˊ�"�W�Ck���.�PGA(aiHt	q�R}I��
Xzp��{�U�~B0W�j�=����8&a��������+L٠D _�$�o�e��=���x�/�}���aT�ot�.9k���};{0��Vvil�~�yl�el�ے�ԫ�W�]��q�#d+O��z�D�[�ڿV�:�r�(p��>�� ��9��͞�j�kZ��m��!0���]�M�?���*�,`aT�˘7E'
���4*����"����yqlE����%
�Y= wh����98�S��y*!��%͊S�����:"'��;�^ʭ�5!P��?��`%��KOӯ�.��]�x/#��z��O�c��S�{���=5�Þ��<�>���U~`��>�$�%	�<�p��q|��J{��YH6�J�1�tU��ِ�Z��h���Q̫���W<���PI�V
0q+��*mIV(tL �S��d��/;��N��d`�;����1 ���\�/��q�4�p�G�N.X�aOF p��I��Kt���𜭵���@<�S�g���� �sX���*a-(H-='m����R�6),$�&�G���mc�3A 8vA��Ot�3�]�!�j���Дs�s�"H���wV�)$0�JRV|���N�ڔc�-[2`����h; $<v��3�<3�2T
FZ��_����"�b��(�<T^���N�fEͪ"1��\����3<gLy���U�9ՉA������j⎟��H��=���+߮'mmc�7�=v�j���U��s��E�"m����6���[]�Y��؂f�?���zO��ت忱s���$�E���Â鿕 $�h�:I��M ۻ%%��L/��D^N��^T"�gn�Z�yve�����8'�uݟ_���mݟ�gE����!1��ዚ�\�.Ɩ��>aP���t~��^L6[�1����1�&8�u8ӣ�|鹴G�y��}�%;[�Tq��yi0��/ǚ$j�>"�z�>\����3��#�yy��'ℳp����%��Y�z��$u
�%�O��Ѝ��<V���"�çku���KM*	t܇�h�o�����y��fx�d�E8iK��of�����j�:�D�����y|��Gz�N���8MT!��A�&���TY]�x�풎4��e�1����'\Q�眺��/�3���˂�xhTZ���-{fU.�y`i�ZKH��w� ���e�1b��ز	x���6�(��t��ύ�i�Y4�U��Y܊�R6o?��s���/:Qy�%����?�"�%�V���tgW�����G2�_�o�o)f��`���/�86=$��e�"=u�]�"�b��Q�0A�����5��T�{,!Nn�SnZmq����@���� �Y��yi*� Z�Yb�a�E�ď̓�g?A��s��__�V��4�IX�������0Q�����fN��@.�oD���\�RIg��7������M�i7���"b�� ��{�/%�{M���3SW#޶��C���Y�EG��Ǵ+$�|�[�d��a�S�]����Fhg�f��L�L2�5N���$�4��y F����Z�k_�%rٝP��m�6g�VF�=*<������6�Йx����1Zi�䲠�)�M'z�TG��;�|�G�- �
��.B����#�jl����!�A�5���ON��~8+�_��i���:,����Ӿ�1�'�?�⏜�XD𓷌�<1�����v���^xH(���P���2_���Gl��.6�����fؤbp��	�4�x��M~-)[}촕����!�"�Z�� ����ǀ����G ί�,~l����%5�D}t�!7˵2 ���(�O����t�a�r
��,��4T5��SA���r�xep�5�pk�&���E���L�E	���Q���Lu�}�^���;�^>2�f�Oo�L3�~�k��f�pv����Ho��vH�u1)T
�uB�x5|'fH\�ȨVIV��_o�Lz�#>�v.vx
v^�8�����
������?I용��q�΃&��3KcPWR==65`Z��j�k}~�"����B��x�"-�W��/9'8[���B!����X�t>���YO��e�tC�P�,���nPԽ����#9M@��0�)MH|�>�{���Ū�4�OzT����}2m5��r��5S��k�QU=~c�����I]vq�("�������s�7���f�`9�XD�\��:`��ņJ�)��_��" l&�dd��*������� Do
��o�UKl�ղ0��w�8gv�o!����P��� {	G�.�8#E�xm)��#�r��#Ao�tX7\c�6�'�/Q�*�Z&g�~��q�믖�!j���7�n�ㄞ�} �J���������{��M�:5���˅ x#���V7K������v�����z����Պ��<���s�W"+�B�'}��.[�ԑ�$�`����M��P-�r�\���C�?�v�&[{tB~��:�w���{Q*	������7j�9���w�ͻ�q�1G�������~����^.�ġ$"���D�����m�6��Q�ۢ����uT6�[���4��ݙbC~���q��h�sS��y��G�Su(�R
��z�ԭ0h�{����,J��+p�l�pK=
�f+|��x�Ӿ&]�Kn�̹G�0��zYd��!߻��ʔ�N׶CP=���@N�5�d���y�����l�w�h65��+EWQ�n�rJ�/U[���LB퐆����E_jN�&�(���%o=���/�J�qe���.-�Z���QUk���޶��o�U�k҇G�*�u��,�j����z0}�8�	���(@��(�������\*���u[~��h��R��k���Ӣ��|Du0���"W�7I�!�e�Q^��U��k��<���)�����l����=o��;��I؅c^����v��q��޸�g����~�U_I���_���d����n:��}������ �!���#廘Z��0�\��!�P�2m�B%��"�МT$� 0��S�vrpJe,C@��4�y������5�sOi#ϲ�G��TQ�G����vQI���+�̳���L\�?��K��"��c>��Jd�<���
A��t�94>bY���j�U}_<�������%��o�ڤ5����m�*���
+����X�S����Jg�m�� �m�#~At}y��XEgÝ�q�n�[\I���̀
V��c�YVmji�%�8Ϗ&	�t8�w��������Q1��̜����I���>� �|���/S���m���8�,����t��˯,E�} d��i�F%'n����_��D�TpW�aʊ�'�X���C��]Q��C0���CA��y�<��@{���qW�����?��нS��)����Ҟ!yp}������.�_~^u����F?g6��p���~�|n��/$����0h:�׺N�EG�ݏdvUL�#��u�����FnSH1i��"j��� �|z4���(��ͧ30����g@���ۗ�399\|0ƿ-�"��Ҝ��>;���ci����)�g[z	��h��j�ˮ�b����?���ÁH<@-�Ӊ�X�|-n�T��kP��VL�m�$��*˙$���m� �tu�H��A��3GC�I��~����qO`Ëk�9%D����A���[ǖ����W�0|��/p#T+�PIj���m*�9<ί��J�S{f.�����;�츧��`4(>YƎ�f'�`�;�����J�����%&
`�'�;t,�K��a�;��G�t�~�զ����492�@~��-<�	L����-�L���o�2%Si!�.,z,6�_}z�HYj����H{t����z3;�C� �����~���6F�;��<i�Z�s�(C����[H�u�ԝ���㛫�,��X.(�-��~�ک�j�H{Pn�4�s�L��q`��22L���H��7 {`�}��'
u7���j��&*�9�)f���n9.L��B�)�,�szԜ��yJXjB���qю�RU��k��	����M�_,��ݚO*��WJ
��Ȫ`f�.��n��	8��t����@C�(ŀ19���d�<����sd��n��Jc0c�E���8*������ 2c֍r�[�����'so�֪�\�BnO�>�
yŏD���t�Ђ%T"���P(��{����eZ�_�>/=�qȍ-P�6��Й��@ɰܿm��U$�Z�a%Y%�R��k�8Q�@�_�3��4�[R�N�GB���Q~C��Za���uC?��;�$�̆0�%�ڌ9Ol �AnM׃������Q����,��L�|�)��ncɨ��CF����L-�z�(i��z���hR!�zŲ�����Q=m�(Λ!��nT��=|�ڕc=&8�ָH��R�ўD��O��x^iu���J%K<�.T���������N�3�b�
�I�ƶ�G/���	"��.xuR�;򻦌`����y�X����h���Ŏ �6��J�l��5x�Y�#O�E��
��Mf��3�oy}�QNƱ���6���!/��+S���f���դc��%X��]aJq�U�xd������&m����u�/i*�#ǿ���T��$Ҍ�.t��c���٩h�ޗ���Y3�|G��[�h�
���<uPhDwB����:��1F}�s@���H|��6 S��j_15}��R�ǚ�t��^5�l�B�I#�Fm�>�ڦ�uFm�B�M�X�ݾ�J/�[�]�7?�itī�����7އ�����������UA�$j����;����ctjI�u�CD?3""Ye�Gr�5[�~���̑Ȇ�Z�R-Y�1�=�#.�RF���ڌ�E�u"�["���'%���� i&�R����2P
�.�}��@~���ԝ8T�ӹU!My^��!������)�������$j�;��]��+ص!X���g��i�,�� ���{l}G5�Fu���F���ߠ�����9��@Ǝ����c� >���~B4��#��II�= ��3u[��& ���yr�YÙ���p�.�]v��F��X�@���aRe�s�{���w� r3+_C��fJB�h�J+��Jh���!5ɝ�I�����x�p�f.�Y-b��4��D�����c�P_n;�V)Y�w�� �`3
ռwz���$��������Uѵ*>�	�Z�(IٟA�U9�}=��k�:��9����(��4�:�>
vub(�`���O��ܹ�� ߩ2	*�T#F6��m΋��
�Ow��쏿�@��D��#p=j�Ι�[̖9E���W�
qy�KC�$ρ��7r� (#�z�P���C-k�pj�������fr=�C�S�F[+����i��ld7`p 0���P�g�BV�:úT�z����!|�sUjm�x�	��㬘�(�Gr��
y�\G�U��O��Sz���ԭ�}�p�u8�ꏆ}�/�>Ob�	�!�d�QS㩓F�Cv1_w���L�,k�4�bJr �U�y�㥄���ܕZ
{�{༇pb���I�`_@O��sXx���ܗ����8��/$�;�ԺwS3�ۇ��g��.qޞ��0�T�Z�9R�|쥁Zb�5�zpa�{��j�8���P"ݥrd<�}ȱ����pCxjN�3�2�u��C�N�qo����C��o������m~z��%h-���]<-&�� E)ES�]���P����(�8���L���M(x+�����K�v��ֽ��u�e�\�phy��|��|�Z8}��;I`��f�`�/)�џ}����VMY�WlI����a ��p��i�u)��K����hx��r8-u,Bh1:x��K8�&�YI����m�{<�	�H��s] �H���}��V�WkG����U
��	���E	�!۫��bV$m#p
Ɓ��cW�PB �3��F�â�6�4���)I�nEڳ��cs;��t㒼�!qnפ���	�%on��7b���J,I�sԲ��I���}�!�E;c+��(1T�d�5fJr\�8/?�/!������&�[Ɋ�X&X�iݞ�)�$��+�d��/�k�%8��/���7+��]��v���J�l���`��a��Y��^�n�㦏��9�pn�gU���ꘒ�0�ЃV�E�Wr��:}b!��-�N�v\�:\�u���B]XC���Z	�i۫*@|�c�m�P��*'�L<��W�(�U���A�u;t�<����%���!��>nnH�9�+_��砙���fBM5r`�0��]��83�{J{�H��@�lؚ!7��ک$͵o�����P.-��5#k�'�z�wG��{��8Ñ�!+��R���(��>+2'i<5gƷc�ħ&�9;�3�x4=�/<��K<.���zD:��G-���u��̶�a&n�R����T:�p$7Ç��¸E&�O[��d�A���C���c���׃.�`�T	d�{e# $���v|�ApAD,UV!�A�聟��G�"�Ko�'Ϡ�w�׽h����!&����g���*�C���V��Ih�mӎ�X'�Ϟ$T�1����p$����g:yT�}jx+��680�+6_Ok�q���Z��54ŧ�  b�Wu+�X�PhuǸEY�o��{���>����!�}�X<|޷!����cu�������@M>�uJe��j��P&>�c�͝Y׎v��=��Pŧ}?��q_����E�~�=Y�>>��=� �k�O���Q�j!���PY��"
�|�]Y��v����ݜ$�5<x��2����{��νஷ ��dc%[�̹�8t�����z��!�z�r��?���0���4�J\��)�w1%Ӹ���v�hJE�~]��H}�7��P�9�*�9��e`���:�>������G\��P'56V��r�,�0�K+b�L#3��L�*[ �:
v�@��%o����[����=f��q��b�L���]a+��lm���w�_���I(�Vݡ������݄���ʺARF��ul�+��\�H�M�D���y��3�za�3�6EoS�G� |$��)¸�Юz�#i"��y�+}�&��%���F�p�	\L��i�G�^d�ݶ7mR�s#�M&���o���+�P�AO}3��N��,`Z�653g#�x����2����.�l<HRO�'��*��x�]�ٸ���hy��oɴ�ȹB��U�u|ivף�����\���ɦ@��=Z��%����C�K��At���/o~[f��c�(��e��al�!q۳��v��1V��K�|G ����pK��e\��mV��lǜh)w}�	i?��̙܅�B�w�v��"¾�9�,��������U)���u�@Ӓ�����5j3�0�9��p�M�F��tب��Ft����&7�NF�"m4�M�K�ds�/E!qPn�Ӻ/�\#�n��rPrG1��{����6�Kw'H��n�s-�luA��5$V���%��@� ���w����S�!�P!��ܭe�B�,�=Ư���M����j�P7��Ve�z)y���,J��o*Y��F���1M'^環�!�ZP�aq��I;�?����e�UZ���pGqt�dR��j{;؟f��j���
GH9{��$6#��ͼ�IԻ��t���%>jq�4]j�?X�3{�?<��[m���W�r�Ѩ�)�sצ�Wv�����߿P^ڮ<�aؗ>N�BjYd^yW�l[4j��!lVxMCOy� c�l!��aA%�P�t�G����3E����NRԦ��J�'w���2�d�!Y�t�3�yBlc�vs����ȵ��F�dk/�ґ��4d3�d�!c:2�ͨN�-1�l������&dg��m�����V-���5�Չ�ېG�ߒ�����F|�R@�7҆��<��1�Z����ۖ��j���.��f���\̋곹��%~(������x�#�C�`�e�]�V�0�(COD&&�r�-����m�?s�:��FP��
nP"���ƨW��J�d�.3���H��\Sy-���ŉz���}���P?����o\����0��&���{�Dy���jѧo����]�v�:,���
��7�`�N�6@F�{h���Kg����MG���{��Qc�&[�Jm�쿾���b��%�pA�ODa轤y�_ʪq<6JN�P	.�0��ke\G�ڕZ�=�2�yx��cct�p�)��գ��hi1��T��������ڇ���<����{m�U���?�W�\ ��5k��L�����
;K����&7��d%%�����:C6Cz=��#U���2'���ڞ�J�k�s�c���?¹4[?���p/����@����w碌~=JV�6=��)�Rl�u�z�_���5sU����� �QlO뢎�ț�B!Z����4U�U�2-����z��2��Ve��t��q ��H���)���+'c�l{F/evH`qz���
W�KG��d��l+��B.ּ=�k�<�����҃D����f8�v���@ػ�'=���¬\���1J�2ApSB��MF��H( ��!���N�b������}�c�A��j-{{։��.)X����t���L4����a2�&��C�#~����e5�fS��I�R�8�����*��,R׾-X�������&܊ʧꪵd�L��({���`"m�j�
sH
�+Lm��
v�4����pp?�4)�B�N�2>��pR5&�k��Oz	�?��~���{�hYN��C���$e0n�=��ـ�<H���K޶�&@2P}�%#�Rn�An��ȕk�SGް
ɩ���qO�wIx�ٚ��}�Q��g�{B���ܖ��X@E=���DK&��� �C���|L�^��"J���a�K[W?�d���iNw�~����J�
Wq�����%E���L�1!�"Œ���_�����j�	,+�}Hp	�'(`s���)g�D��%R&s!A�5�,O.�)�uD*X�7I� �
��C�zx+�s#
����V�QM�������?xP�.EQ�Xl�x����Q["ǎ�S�����.���A|8�9��CR�P��*�۰l�]J<#�
LP�c�8��ҩ:H¹��86,���RQ��X]���IA�S�~��nn�㿇��²���Q@��}_{�S�uB������z��5<V��z/o$g"y��LR��Q6�����+� ���5��[���m�v�QS�*D��JtL�A������� ��>ZMS�.&}��P�����B+;��i%��w����>��E��A}��r0�CI5,��:��y�^-�*�#���W��nʌ+�#VՎ2.��r���5���Sq-%[hmp�p��A-�(�`�th@��n�;�:����y�s�؅z#���iX��CJ;��d���!,�������-���+^���Q�T̍U��Q�뫺��ζJ�>i�P����A�h��Eg�-2,Ԓl@�x�9$�
�O�Jss1� g݈���V�R�{����C�;�G)�ܲ��Y��U��EY��
7�`�]cS¿ˆ7�O3�Tj���D䢯�k�[X2�偗��g�d=����o��)������du�%�K���y�8�a�?uEz�#e�S�;DV�<�톘�貀mk�a3�	�e��������d�����7jz�����]f�Eq�m���8���n �o��f��w@d5���^���!w8�t�Mf7�Q��p����d��5��q���xp`�/f�<tI24���C���8D��~�y�K�� �J�M����,]�'h���S�B��r�+���	ݍ����P1�фb�*��9r
b#�Ay]ߏa�?�k0^�v�����5�ȟT��}�h��u�����a�;Y�t��rIp���:hyE�h0�v��[M�ȑ���B�hS�b��D�I��^v[%��R��Tp�E�9Z�)Q{�(hR������J@U��NN!�j@Aq�L������.V0"�!�򃺏_�u�]�5���,�r_�����3��t�t��7p,WjVkT�{�u!QY{6{9��B��z��v�������O�e���ٝ�R������
m.�!�lq�w��Uؤ{�bR�už1z��d�,�����+u�����ȼ!ҏ���v�g�Y<��������~U9���x9���S�#��3�s�6��'=Ӄ�z^����YX�����%�ZX[vZ|�7���d7�y�݃!}e�:�8+vx���F���u+�S+�U�����a�x��5��Mn�<K�bk~W.%����3I6�������������5�P<Lߜ&��a�����h�"������Fݘt!7{y?����T���ɥY��x��}x'6��p��=�"	L��;�r�(����_�-4�V[,[�.�m�/�H�b�"E��٧�����:W��ȏ'en=QBV���}u����v�
��"(AUm�K���GCY�**/�U�u���B�ө�,���6S{��&Ӣ�du+x+1����u߆�G=�8kF>ʴ4����/�#f���3���$u:��x��~�+�y��,u��=�}��
e��W�>6Y݆+��M�%���oqs�l%�g�2F��������3E��E=p?}�S�>�SjI�M5B�6�7+�zj'�.lٷ@��R��Cd:�7m.�s��#XK����,�p}[�����&zT�a_��S%`�	�'7��[��#�]��p���M�)������!Q���V:­3'֖.�d��k>�r�L�x��w��( N#�U<��:��Jg�������^��}�~��u�p���7�n���r����֤���x��y����+º��ܚ�럭�뤐~��+.Q7q�PUSt��H��D�O"Qcex�V�0�N��F$���n&�/Ѝ�\��C�?����m�^���7���(CF�D�����F�u.O��a�KC��!In��R�����oK�)=l0�
r��Iv��z0��.���0�s8�>w�������@�+&�j���Du�ԭ]�a"�jy�D����ׅ*�x�ؑ��* ����F?<p�,S�����g-"	�)S��V;V0�1ʈ❼J�i�2��%ݗz��e`�t�����O:�d��\� �Bw��s��s�#������s\
r�;� ��?hQ��Lc}�ϟE����X��e���u�hg�P/ �i��a4�F �w �q+���֢\4��ؕ���wY�"=3��z��1F�4W<�<�v�e��䪊�-==�/
�@{��_:$]l���@3�ni܉-��K&���cFp}��^^�h�wbH�d���y�#�ЃEɵ�u�+�e�;�?����T@�]*��@;=|>9�
2E�#+��6����DP����u93*W���fqߩx�,V�n����W��Ι���J#O)�_��|�[������0 ��"R���^�[8�����>�����l�?�]
�hmA
��#�-��1�f��2c�[@�^�l��ᒤ9P��b1�8�����*��Z�aUA�S�l���&e�V�·�i�$�p��}_��i��kX��g��ˮM��F����a��u�3q�;����*n���hf�إx�9�������X�vo2�#�u������V��]/��k[1*֫3�w�.J?��&V�:~=i¬y+-�5z<y�0ao��d�|�������{�҂t�'�j���[�MLQXp9�� p�w9����*}��X�^ ��)�1yF�A� �O8?��ꀷgYV���b�D	���d�o��߀v���-oT����á�GJ�~�^�����d�fa��e��w�F�Z�3�Z��)i��:m���1��RPp�ѐN��3���iP믞v�]z���Tr\�}�����S���l������ȓ��bc��Cv7�2�}������.,�`��S������y��h����-�i��(D��H�NU���Y�~��ɢ��C{�^u6!(,sA��f艾�Õ�se�m��NL�i\{�~>��;��9U�^��Z�^Y���]}&�_h8s��s��		�;QNҥX�6�q*�$,�L�+�:Zg"����7��h���h�4,��Sq�R/�鴖��@�@j�E	�4b�����$q��z�?���G|��D��(�u�?���w��G�lvRw�z��a.�5�������b���W�l����3�aU3"!|�=g��)��]{�^��y����{c/�?yG���ټU`eD�wR��D���31&�l'� �:�?T��~]%��=1���|�לϖ��4�-��P����}v-g���[�u�QC���
���E�>y���8@�&F ?xU��4w0�$HC�x5��e�z���qDH�����\?��>2�ٚ��Fƃ�S�{�}lm���H6���l/���XK��<��!c$r5��թ�h�I���w��Y�K��LZGJ��UB�&�����j���g$�[�HL�?��YneLrl
b��[��o��f	�7<�5��|�mg=�wh���/JZ���%r�ow5���N�=	F�4b�uS��m��/��z�j`@�
�˾�p'b��*�C9��{��ĉI�8>�.�ʜ���.n��'w����~�z��0?�&H�=��o��w�a�p��!�сWH��Dv�0G}�o�Y�$�.�҄���z�E��$���f���w�;����A����*e�3�
,��Y�')�Rq���w�xGK)�S	���T;Е�Z�$���4�-֠�So,�����_�h�����vp
���{�f@wl9�2~C2r���i�� �	��k�D�龎̧��M*�u�ݥ��D��a�S"�Jc��Y��8��<��iWg:)��-�U�&x�ַ/��x8�6
yG*$-=���/Պ�^�0��W�C�� ���\�M�����U��)7����N������w�b'�:w2�c:٪�z}e���7!|��l�1�w�!e,�**?4���"�|t��߻��cjJ8(g�D}�vj�H����kkCi�����L2t����)� ���r�VhP]��P?� ��%о'�%���F3����gN���ok�,�{D��<���c�I����u#��р���
�L`�L)N���GD�D��[�K�N���\йN7[�b�Ӭ���7��k<Py����kIk��@�� ��#5rFD r�n�Ŷvȴ<�Ѭ�V�Y��fݸa;��tv�I���$) i�w�l/<f<Y�<b��4����h�o��(����<�1,��N;�TV�8�pS�:���~C(bJ+8A����t#q��$�lj�TZ"*��(?|���Ṉ���}��+9�c�rh�4 6*�{��S;Mؓ��ZW:$�ά�H��l��:�����>����UDeUas7;٤ڮ�I!���������<��gP�H���2�/�z���r)�qǰ�#qW�V��aP��&]���1�w��~��һĠ S���%��N
� �E�Be����o��Оd���t�ba�2	>9h�(G\��P)���UsQq��3�J�M��X�v`�9�k?�z?~K���3��M; �_��ph�eU�����7��yr_����a�e/uQ�N�C������n;�cE�o�疐ZU�BX���BQR3�[������q��eC��% #b?�����I����6�ʶ� Bl�X��y��,���ğ����3S�>>�A���~~ ���<v���v;�#��d�`��#�7[��-Ҙf-H��"�蹠����������])��<��ۻF�$��4깣��&�����܍��Ų� �����G^�{�Xrj@Et'�Ķ��Ø#�q��Z�cD� B(vά@F�|��q��k�e�l���k���gx���Z~�6�OJ�d&8����\�3�iK�5�E�6y���B ���e�X��+�x^?��.��N�Eg�~}��s�XQQ@��>KqG覾�o��z|���a9��5�ޤ�S�<H�K�0�9���"�窎�XD��mՅ-�~t =@���[����ᅣ��m庪��<���������v<������I�x�/<#�s��g��*seR�	�.�DX�>��G�r�9��.Mʭ�e�!����ɤ�E\!V��O��ʇ�J�a5;��{�����0����ټ�QUQ)�
�	Pq����,���S���&	k+�zBZ[�7t�c�0K˥�[<bp��B�2�Q;�DE����ſ�\D�5vu�A挘�/>���f�(iW�yz@ͪf�}{���1��A"�UU`�<I'����j�혨>m90�Tܐ�Y��\���Ā��*��-'G]kv1oUt=���lլ��
�;8�pid�|�����褌`����|���������"��n(m�4��*�vP)���|"�IL+N��ʥ����?�ԫ�R��zID�[H+pd��uA2x��80|z��?a6���{�s!4��?9z��^�ۀM�!�RL}'Wd����4p�&�WW��R�l�E�D�O�ê�^�^��W	S4��㔕cm��.�+���EJ�d
��W�TL<���S�k�o15F
)��s�!�m&Vi��6�kx��O���}��L�A�@��븪ڹX:d)���WC*�(|A�h��0�TۯWC�}>���
��Tj.����3�^HHֲ\`�{Mpnp����?����ʰ�G�σ�ٕ�k$�:o��j���|+Eo�K*��\�_r�eU\�a�U.D���Q�9	i��}��X�:��hz�pi���$&+�cS��IU4|w�:_�Ɯ�P��� ���puÃE��:�����95h0CW/�.���WK"�d�O�Ob��5R�2ِ�/���mI8��{Y�i΂ɽi�t���ی�o�d<�T�ps��"p��b[��sU[����|��_�����.č�WF������wk���,�x�~�ܩ�}��A�O��-%�O�6`*DǸ��i5=�Fb�5�4���i|��lD4�@>HVx`EfHn*F\�~:I�CM :�wDz�j�O���<�;l�S
�=8z :& Il�}��f2=���/�x@3��ZUف�N�2r���%�p���ݼM�������R
�D�<&����5?��JW����w�������E'�<vB�x~Mt�5|�����xa]'��a&��Y��*l�$وr&�D���I��!:?�� �3`Mp���;��B�.�kV�j�-'l��VBS�A}DePa�4=.K��Hܿę�*��@��r�52m�~��\��B���#�4S{��+>�1��wǗ�rE���N7�w�qmU$�K�	$��	�ȝ�]��N�pR�����"�$�r \˩�iN�qu����b�c!,�C�5i�x��n=l���*�	��v�Ȍ��vl�"���J0s
��?C��k�B=l<�&f��07w#�v�i��q//'W4PW��(��(9x������Pٰ����u��6����!�v�+����P����<��f�C �~��.H�!��mf�-��G�&y��������=�_FU�:�2. X|�>a�����n�t	�"d�{�mG6߯� U{&6���/e�h]���ꈋ�{t@��:Q�����=�"��..I�X<ɼ5���:�ot}��PH�F�F)c�y���p����p��Y�� ����c_����帟7��͕LS�:��H^�w4��9���l՘d���|�p�FkZj"�5(�Q���z�p�c�(K�~s"���v�pȟ��f�JL�)��q�T��z|��*�T�q��~e�&�v�W�O��Gd�z�OUZ��<y���Eݸ�;@���߉�`kH�����Q� $�L�J	���٦�K8ڻ��/��w��}q�x��5��� �pqGϩT�#���� ���l�>����َ}�E'j3h��P���`�ѝ=W8[�{+Jy�F��A��'��!r������\|��s%ִ�S����Y������`���=�T�š2�Ǌ���'����B
nQB&y�ܒs�bt_q�]�[�ϱ=m`���/�����H��`��u1���>�ycn�s�ɮ�^�C����`��_�䒰���:):K���"ίJT!n�e8��ҷâ�8Z	�>��ݲ�9n��Qf��hJ8L8�Z6�UwZv�3�� e�+*�/E�m���tm�y�������lQ��B��w�Y�^Z
�v�#�A�3��ݎ-zc,�z��$��& �u}8\IRn?������]��s?�:L�#�����q�(��(s�L( �0N����>k�]�m�����D��_<���u���t/E��Z6_�7<��gߔ)���]��T����ɌP��sţ8�����1���!4���Wmm��6��-�$HWj�ܼ���&�`$�yO�_�����}��{�*\�g>�R�{����6�c- 6���Mޚ����L�Ł���|�Q��
���e"!�m��-�;�K=R���� tj�Q��Ո/Lߍ��]�5`���Rw	��J��\��Lp!�?yʋU�"�/O�lş��q�כMWQOު�ud�����<+�a��L�`�R�G�	���n�A��SRVT�	lo4CH���vo(�}�qA��^�/RӐa$�+���3
�7ס����յ��O���>:�].����t�[~ҙ�2�(�����m��!��;j%.�zƋ���S�xt��y��Hi�ޒu�̔"\�O�����|�܋��9�Y@2��U���Ĵ���1����l�,	'� 8�X�#A&��Ih��ۆ���֒�2oxa�����>f7W��S��f�;�nb�f�����t�R^GB �M��.�BQ]���@�+�۽�F/���R�����i�0l�;����M�R;|����;��*e����0�Yo������YU�2��b���^7휧�\_�ȋY�>���u%ݒ��5X�T�c��/pZ�=~TuE��0+- ۮ�E�Ai�j�|��dS���w���t4�ud(���8i��8����b�՘!�P|J�@�Y���oQ\r/��Z���˾�^ 5�� ����$Ϯ��-�r�K�U�c��]2ߊ���2�� 
��;��.�A*)��c�tY
u�X#�vY�Z���Il7>��U#��!j�H��v�?#����	5>S���yj3�U�fy{6�#)-�p �ʉb�W�E�Q�<��n]�.!���T|���։#r/Xk����-�B�!Q�A�$hxN�ˍi��_ݛ@�uB�(�[ѹ=��+�k��h�J[�e�G��<��+p$��e�o����ħ�+B_�4�׭45v�5���x�*��3+���b2B����P�~	5�CW�մ�o�ԧMj5g ��N�s)Ƽ `��++�(�*�n��59�c�)��E?�:w%s<���je5�_S<�@ܤ��bˉ�����&���C�F�-�!j�!�y�N�k�P�N�Tד�
�@\x#b#�EU߱C�1����΄�����y�y'��IԜ�+���`��i�7F���q�	��i�������=�?.%jL��W�@��fbs C����k�ڂ]��<΂"i�C~�{�:B�3� �dkHT7�ì�N/��k��ȧTg;1`{s*Õ�q�9�V����$�2���J43/��@��\`�rO�`c'���
�1���g@�k�s^+n��"��2/�9k`#�Ok�ɸ<���2e���1������	 �i�<~�"�M-�����1���c�yN�-?ɗٗ���Jj�T� 1c�}�8�s�K�Ӎd�:��b܆Ȋv?x1������дH��| ?h>m7S��\�zH';9��-.�َ���s�(�!^�)Ӻ*��(װ�l�#�mO�s�~k	�"�A���p@k����i�-��^r2T��<�X���U	AyW�:��v[V��@G���R���ۗX�;���w�ڞ�/9C���J]a�r�
�m�T�i���\�)���R�{Z�"\P-c�����0����!��h!������fE٫���a��6N�����{m%}f�d�~���K"�Ү�?�'E�������������ݳ����%�]>`�F��/�2-�tA&<+�洨��U{�uk!�ub	���q�3&Bq�e�QK9oq�|�{�/v�O�s�>|
�{2��s&�P�0���C�c��0�v�#�5U�[�-��Y�B�j�)���5���Po�r;l��Zm�؇���e��� ����zc)�}S�ׁ1Ri�0��k0�\��##��cf�-
�<���T���߶p����'�k�딜��5�pC����{��P�9��h����eQ@R���b�R�#p�
I9��f�x\�����aR�H��W	�����F�8W��~�D%xZԴ_S��X�\��p�PѮ#�����Ds��3߃�����uB.�
úDʾ\�> �����p�����Uo�i�ۺ�S"�	}�쟻�0�D��x��u�0Z�0���ce/�v�?=� )������r��őB0������h��B�4Mi-�����\�U������Ks�O�&0J��������3Ă���IJ٣Ʌ���sl��O����x��7V-k���M��5Iv(�E^ke�y�%������R޸���� �Q�\�\Pp����*8pa�:���>��O�9�%�Km��=S.�&�%S-�mϲGZ;R���������+P��Us1.�'�#��b����:����������F�����W��?�l�������d�����Ѭd�CU���V�/a�	�k��*�ta��ELݓ_@V����oms�:�x��L�wp8w�J�k$=m��%�a%�(4u���w%%��h��G�>�\����u��]��!ҳ����}�S'���`��{��j�����a��`�N��d���~hl��
c�$-j�A�13��D��8�LM�\��);*T�rBWƱ��0.nW�e	�|�/7�ަL��F��:�l�|�/P'��������!��:���{����C=��@n���/�t'ڈ�롺��_�{��[��*�7W ʹP�ZAuByt����T��ah���#-"֦J�p��Q�V8�u
��BPY�#P���,��*�P(cX��WQ�����=��	J�[tDm}(�N�p?���C�t�Yǡ%N�lFJd����w:J���"��D>��U$@JJ�p�P9�\l�r����t`h�R��֘�t�˶������($<�^���-:e',.�ei2��a�yu��]��i�)q9ebWNg��|�o-5v}��^�B���IR|bw�!�������(w_�j�\7r�,m[f��B��a��/�6g�����4!��1_��@UW�R���_13�D��|=��9/�$n�{��L�i��* �	C���
�v�Ƙ�!'�a�8����?�݃�~�IV.�օ��%a�!����Vaf�d��3�x�j��!K�TתǙH��_�9�ˇ���ɳrP���/%��f=%��>0�v�Oe�2S��d0�\=�Zd
g!�RZ�a�0�%�O�� )���K��I�2!�hT��Ǽ-`FqJ~N�.��0w7o�2އ>k��[��Ww�]t���l���T_"��S.�U����1��������ǌi�M"���R�8����1_N/� �e�q]��w;�4,d�Oh+�f��A���8�e���ę���{kÚ��~r��:Z��������B��(�;$ID��y~
�Ԑ�4��F}J�I���u��K*�a����.N�#���M�)I6�E��7 @�xl���BPލ�婂5��i}X��}��Rb �m`B��0j�B|�;���x��mʙ���Ц�ޓ�`���O�^6��=H 0�|��K�q�&됋�s �	�v�_40Ş>��?�
�n��
-��WQ�`g<�&0A�SL�/��:p����m;ϗL���f�s�`��GN�yƎ����zW�T�*Ps�)Q�i����������� ܍Ӯ�'���.gT���}�z���j=���� �W�곿����=)��ͪ�q��s���r���:?YS������N�?����v{��#��ϧ�3�-Ƒ�l�^Ce�Y����&S��\�ò¤^L4�*��p\x�I �� >�a�5^8>�'�?Q+=� [�k�1�I�7��X%|P� (�y�B�����#a} a^�����x�ns����^+ͧPUE�&�k�Wut���ǣ����{��Zle�Z,r=��T�&�#�UV	ѻC xUk�{��?�:ڄ�%M���VĴ0!�_�45i�Xk_'$��$�� ѣVOrn�츯�p�IT�%��(L��Ϡ(�S���ˏ�[�l�F�mE�K��'��fmZ�";2 �,斌 ?�+��F6��vYxs�f-P��9`����j�pOA�q����D�)IE��S �������bt��)���
�៱����P�LW���7�Ң��^��6g�X���z6a��G6�]�̓YɅ��+֩��g2�]�9�UY�tBR�u��3:_����G^=H!Ϝ~�L.�p���&�r�"�[������[x������H���I�ky�k�ΧS�I�@C'/Xp�u����^��I�n&w6x�a�.@�h�MO�ݹ��`#��w��Ŗ>�9p`r�7��9=��ω�G��k������l�_��G��@����nu��;N`U�W���H������q(G���%�	H�@p#�q��'��w���<�7���G�~��ǞL�cRw��	@�I����o��.��*���L������愼H������tEr<���|9�5+�ӂ�+B9���Lf���|���m���S
vu�9�T�R{8���?�~q��g�^?��o�7<�8;Q�͠��C�a�=T1x�CU��w�(k{��I��~{��̃�?'���	��@�����؝A}��s�M�߮��&�mYy������h#�0���,��R���C�&\
��D�T��I���<���U:�_t�8��A:WQ��4�Oɴ�b_>3���e��dX>?~4�:��c�. �q�n|p���G���Vg���%�`�g`ʷ8@G�q�KZ�ך��/��Js*kd:�
��eC���H����@� *�36S��	������z�mؽ2?ȭ_>ʏ��IV���`jGGn�D�wC�K���w~��t�������K�'�����ֳ��2˚�ՠ"������u��E��{���S�{��&�}l9�.&��Fw����K� ɸ�,�D!n�Ҫ�((�ӌ7o�� ���{�gJY6��ꌚ�G��Z�9�_\):�&]�kM	3|Q�5��5^N&A���|B�_���WO}�p_�b�R�
3��xp�8�f�P���D�Ư�즨=N��|fF��i%`GD ,�ݴ���͗{6��Y7����V�J♝��Z3�M��p������O�k��	�Fgf�U�JTS�q�n�!��Iؔ]��u���_�4i�������R�_]�n���?��W(�i���"
)y�j����k��=g^D���>l^(b{�rsD�!8��, ϕ��N�������aр����QsDQ�%�Q�'�6��M�����Q��T�$C�]�f�cve���F���6�ڣ��&x=� ��K�n��=-���~�k
TC��/�nq��`�H����^��[Q��UQw�̎��|�@}�,ͅ�P�d)��ޱi*�Ѵ� ¾u��{�:k���[F������Qs��VM�`�ڳ�E-)bs�(�6�4��IN4$E�9IҌ�h�ń&��H�cq��د1o���1�
��u�����e�$����j�|)]�b�	:��%�ow�1,|ly�9܂�5BM�b��t��'���[����%�[oH�Wx6�"���_�fy�'^�0���)���a�n:�Tr^��Q��X�ꏧT��Ў[�i���b�j�k�KE�sݾHќ��ƭO�s B����{�o�{l��2I�K����IQ�hX��!YGz�o��p$�����vN�=j�ㄏ�7��
�JPQ���"�E�Q����M��͜��9�٘S�Cm&o=E����Ra54�(��N�fz7Ѝ�XG\bw�T����H��3V���i�|��is�~����;������Ɖn���|N�I��W-hUM�k�� �~�� �1y�iV�5�8�^)�G��`�tHG��w�[��<���ӏ2�NE�������E��V�T$��uoA?�7��gR��io�+��5����h"�I���ggV_s��|�^\�펷t���:��^�s<��/ч2��D�R�����OQ���XvH��]]piO��L�e����j��H�n;={��hζ��::P��q�����9���Lg�<�6k�n'��8�[��.nKOy�1�.�l�3�k�&��x�c�d*l�7S�0�t�
!�v��z��u�$U���)5@��8��!m�����v�� T�O�vh������e:���W�R�C��<J��X�.`B2�p|��*1�zy�R f*3�gD�2���g����y�a�*j�= �9�O�Gs>WԵR������^�D�7P��AŐFR�:�
��H�V�j���ŒO裛��=�S�F��  K̬�Ԣs�p��w�����ò�~��]�(/�F%��H��{l�oq%��X�#�Sg�ү�p������;#n[�\�4Uz��"iQ?�*C_���Jw��G!n�����l�:%�o�QQX�������?�yה �x8mi�
�KZ4�����C�w�ե���I���}��e�Nikx�j�1@������.�`"�|b�8�-vS*�@���j�����|��9[|2��� S��|�o�@N�[KS
�����o��2�4?�?�Js�m�������3��'���%�*��EiQ�h�P8�+'��NFl�=�}?�����ͯղ,�D�rz��B+1aJ2��t��&8%�5�S��e�~�U�F���ߐt���&�E�v�BaX����U	�gY� �ˋ��O_�7�/ �.�Q/�iw9�{��tx��Y�JF��5Q�y�i����Da.4=�j�φ�,�(��r�U�WY�A�l�|�_����Hc�gd;e�Qj�� �+��� �T�[�4	��^��"��e�]�a͸�-ka�L������w�<�����<Lu������S�b!�#��G��}3��積ԸGݝ@mJ��Ln(�D�/Rw��QD�o!r%�hR�s�z �U?!�@�d��b��y��7�N���u���˶(���N��QY�����6�~����ށ�m��j�p+v����g�� ��{2���ܖm�����TGF��k֟�M�7)����Z���9��6ҦHw5�W�Z��6��v=�:T���s�;��PvC�m�d��!4ڹ��|kzI<ٿ�~�AD�{2�6Aղ�	������%����cݞzS�wY�%8H$)�^���=����&�l���Y�lj����&�ۃt�^}5-��̙�c�O���_�7�<�U�ҝ��wge��VZ��ixc`A�b���c�?����kW���שz���N"ǅ2�k��mZ���C��+W�$>{$�zB�:��G��ؾG�X����!L<���덧m�J��7n.�҂������n�+������M�'��	/ϒ�`��R��8� ��d���~�z�98WbA��P[;5�	Ńd�sh$� ��RƸY���L�3����[��VA�^x�KC��/f6z���`%Q����V��;�g����&L~/!v�v�v���@��t��Z>�Y���aU�X�W����������z���;�����߸�rC?6��Ff��5�>E8��q��nNG�k�/b�\2��
�2p;�����ނ缤�y��@V/ǚSf�m� 7�"p�E]&5���e�m�d�߹_�<����@�����.��~(N���8[�K��(��;}���6��ﵘ�n0�x��ݟ�N�v=�ņ�T���3x�B�uSZj2_r�X�φ ��E���~���Zs<���{y�R���[�V`L0O)^#0��˳ŴL��1t2Qً��Ԓ�E��%	���g���v��Of:u�n~;V]�O	�k(`�,s�NZ��B����G��!�2Mi�-�,}'��	���
�iZ 1'�"��@6~G�I��k��xZO�}\�ʎ�D?�׍q��ǉ�;*k��wE���t�᧘��d��5K�;�%��-��b�\���3u�C2�ݼ�iUghr�7C3��e��Jj��cm;��H���K��Y�}�x�5>զY�w2dMbR��C��j��(�1��5��c�S�ۯ�2ǫP4K�<���N�|z�<�증yb�~�|~��խ�S���$�r�+���nt�MH��J��[�9�<��qA����tam����{ß����'�*���iu���T���wq%
��G�u$��?� $�^�0���h�0{�5�� ����3��2p��.>��I����{>z	����G�o�0��!1�y��^�o�.�dQY�O�ߐI61`B���#Hn�%�PRD5#��XS6_�d��i`��H��\�"mXT�e�tܘ�����kR�L�$�2�`,�1*@�چz�@B�s�����,�p�I<�\�f��5"zۃkܷ��&~��Fm���:�" �Kv�v.s\4#��S:��X��0;�ʘމ�S�[_�;��~��W��!�J�,��E^>��'vyU�x�z��_�� *~��FJ��Z�� I<c򋲀���e���]���e�[{\�X��<J���L��,_��VOV�Ͽ��\T��L9&�"��p���G�ZBp�YvA:�?��J�D�����-�ݴ~�y��E��cBn�B7��]���m��cuvq&�ۃ@�+�ɬ]�O�s�,��e�wP���=`�㄀rwt \��0{9�T����$vU㲤��fP�ԇ���}��q����%F���!��T��1-�; ��q5�oeJJ5AXx��o�%c�[p"�!|4�ָ8,�.]�]���-�emA�#m=��8n��Oڍ����~u�Q&���Z�^(�3�@Şݠ�fE����x�EU��J㎻�S�f(Q���'3�k��J�m�	WA��}�3�֤�wV0-.�-�n�VWY��(+I���C�����[��Y`�~���	^��Hs�����p7�%BD�_�z2 Q'�W��^sSF<�����@1�Nl�ݭ�۲Y�?5�A�y ���R����ø��s>S�>)���
]�����<�[�bnZ���͠��=�g�DD}�W��$qr��1��|��;�P"S�,�a���iv}���pO.񍌕���`���|�O�=�#�}'�p�A�$m�}Ka��o&�t~����=���"J�?��{X�WM�����<]���Y���Kv�d����¡����Z��/�[f�Wbwٟ������=�s�YR>�����+3d�^�ޖ� ��_N ��47��=����As�r�{c��8JR���챖��c^�����O����)5��� ��'9���<a�Vh`7=�KzAQh�S]
�.�֤�[�>�{@�L�Do�]��ddTo�Y��/��v�T}A(�b��Yd_��GF�A��b�$�ɋ���&���?��������ڶ�:���WʞJ�,=���#菀�X`���RV�)8��V���C�~�ƥO�����
��KP�ªҒ�k��-s֒$Ώ­�� ���e��n|6��(K���\ �"W��?.�����/�0_¦��n�0��NO�S�+�B����`�#巔�M��QZQ1��~pځ*b���˶k��2+����Mo��r�Y��dX��i��L8`a`͎�B��p�y�	�6��!���s��f�To�����.�;'�Ks��H���;Dc�;ڏc "���򈐳0�,۰�(��.��g�*Ȅe��u�;�_�, ���o��\����Cr?�\���e^�s�.��2;��Q���h!��d�6U���E����_e� �:���-B(�Z�pjt���,�塏�{PT��� �O	���*8�U����Ďv�@�w�lc������ǽ qP�c�0=�#딄:���c:�A(s����4 �eZ��k8H�Jẑ�<<ܥ`R-b�{����m�sm�&)qg&5q*_&�e�ŵ��X���>�D�J�T�)��:JNo��@/dvۓ�[\X� �;�����@�P�w92TA�n\f���6��+�z:%����vޓ�#�#�N���B��q����e�\���H�
1���3$���n�nU̎vL�D��7�;����:M���;6��I�������dt����l&,3��Y�ҧ�]M���}�&d�MV��$�M�0:����H����j� E�����F��=���V�
�@���/SJ���ÆV���c�M���YU�����	z�)}|�;��q7�hd K�b3Q��Po��r�(D8���Qy�>Z��̒\�޺F�8Q��<�A�D�6�}��dM٠X~쬠�aP�yR䒉�F��?5Zd��0�pL�*�H���Y��&q�%B��2�5�?haz���vj��L��d�<:ep;L5��=!^��9�����Ա�1\�m,Ҽ�[p�m�5��0�n�^�ҫWS�6����D��NV{�v�h���K@"���+�!�nT���=�S��!%�����Pj��?	��>�%ᮝ������y��	B!D���`���mr�u������܁��ߗ㽃>
,� æG�8�	Sۅ�{/U�R�l���3��\Ү���t�r}j�籄���� �#�*>��P�"c7��� �����0��)ϑ�M&�vH���A�WUig����̐et��X��$��5��[|�R�o�Hn��J*��d��S+�Օ��+o��ZxCԔp���ul���I��:Gj�"���Q�gZ`��k�D�N݃O��G�V(�!�"�>���|�gqBqd4����0`�?'s��4�`Nf�;u/�j6/�j�P�QG�G�k}�0�:��F%B��`݆�c�֒|����D���ڔ��9��w�l[�M�ģ(n巸5��H��i�	yC�����d:#���������y����V�(?��\#��+�S�j��v,J?����xBn�]��$��α�l �~+�mh-��捓?�5��KbBn�U��mg&C8cf����xh�9�Y����֐A!�S�w���YZ�~Hڠd2��<�hwD	W|������hpE�V���`�TL�	I$.�V!LP{�/���"��M������k�מ��7�����X!�CU�H� �b*k��wT
�����%eӵ3%�1�o9�0�C��f�&�� ���ڱ A�O��{���ϖ�g4A,�lQ��R!+�� ��d�b�Nr�C^/E�A'�O>�8�38��6����)Y|
�)�R��Z0=Nn2M[�n)$�گ��zy�-4F��[�4��U��42�J���Z�a�U�SB�O�L���a��d��BO亊ΐ=}J��qR�5�#���'�����]� �:�8>�O�J�^H3.�A���Bo����(~j)��<kz!]�+�QO��D_�d�������C%�;��S�f�ݏ�Z��yA#�<K�^��ā�+߽��Zt)�J���a�9� ��ፊ���u��uӶ��z,n�(s�SOZ�}E0v�y�l���I�[��;���p0�Ѱt�� FĠ�?���1w��z�,<t���a�`?�՛�����^�'������),�C_���G��{盝��WDpRD�'�+��
��#爍{rR%L5`��F�@x�h|�;����8����L�n�K���Ҫ�(zO'�']��}�`Ď��	ƣ���
yt?�/�!��]��q �p���t/�ڲ���*4)B�#�Qiʕ]D�#�ɾ轛H�Q�r�y���e��gB���;c7�Adʴ����!.8��������dĚD�lr��(�z�� D����tW�ˠ��&�Ny[*��amc�����l����	���t�hF���3j�od��AT��C~�IL8���=3��]����R��b�5H�E� �^P��,Zy.����U�i�2���F����;�Ѣ�-�CD��w��ݽ%bnj��@"��F�C&��=�>�{6 Ȕ��=_�E�c�a^N��ʾ�{��rro5����K��6���n�l4.�&�������2Y��B��ܛ��U�oѥ����M���g��u3͞����h����)؛�*�a?{�jK5[�:H�.����y�^����ʱc��?�QH��hw��{*��3,{���t���|kBm�f!o�.�W��/�)Q�8F�i	جb�|"�����H����M���_���Dk;u�yn��V1*o��_W�̫��&�+M��N�<s��C�����nJ�/T����-�g�}k8�Z��T>;H9=�,'��iA����z�w���^����6�Y�Ơ�K/�6LaD������r��"�u>2����/T��ع%&�i���h�
�^&�辑�"���նB �<�G>8�7[��w����0N*�K��"�������s�������.&��yH�i=��p��']v��b�|��bț�ۓL#�O�?]��p{��Z@��H��؏n��:+��29n����0�3�($>U8�Y��d���|��<��|l[����b񙝅^��a^�%��q/�v����aR�1��p��^+��jboZ�''k��W�	�;��j�Z�#�Mw��֓?~#��P���|���j�&M�S<�O���?z?��p9`y8���ci�P念��g����n �K���n� ,�!|�p������8�A��a	���,���.�� { ^�b�>��M�l�Ŋ�}���H,2���RЇ�]�ص�>Whjq<�AҢCj�py16�������%y?1PiF��K^#[t�"�mܯ2�ꩆŀ���a�_���a���]�[G��+ ��5�)�t�ei��/��q�%���Ǥ�v��.�p��R�EaB�zP����*�Q!o�}������נhm�Ɠ?���;�j�g�}���&ݠ<G��~�����2 '`�+�I2�U�$�5%]�#�h�k�ͧ)c5JU~�Q��11��m�]j�U��+~6 $��v�L�-�Λ
��N>�s�̚b��X���g���ej�o���&L]�Em�9���U�p�|pB����5M��H�(�4��qi��>�	'�Ȑ�0�����׭���>�r\n���h��(��3��|ޯ+�.]I��@N��{7|�G����@'�7 ۛ��0ј��Tq|�S��|�,����դ
�%����j�c��" �f>�.Se�Da�|�Ky����/�]�>�mø�~�Pf��GCY�OUY����e<t=��`������z��� y�ˡ���t���МX`@oFQq�/Խ�w�T�y���U]KPp����`�˩�SϊJB#ff�pk�KQ{u�R���EHIE1*'FBx� ��x\6�x�:^H&�XO�bұg�����Is�٪Xfo�lÈF����$��H�N�y����?6ެI��ޙ����w���@w4gUJ���"oy�`�y�����K|x�\�����A��^fc���	L>F9(����i����{��c���M|v�	饻���" 4�v�����8�S��M����r�%�n�88��3)o�l@��� *.�v���U_,��y���i�Gl��������s�wh�*��l�Q��9����_���d
o9yҔ^����7Ń��>{f4m'
2�9�&�D#%Jf4����g��9���P��g�⩲6������5�K���"Z{`����6��cyگ�΂�i]��[H���RR��wFN
��'��o-&�i�1:*;�uS�}��H��-�QEP�1ՀTfK��/�;���[�o���B1%]IfPbz;'�/[���FhǺ�@��uq���"(�֣�������$���bG~\i�pr�]v�ߴ��n�4�>�'4��
�/���n5��ZʗHO�5��UZ.sU+�*�,2��f>���p!TK_ dg�j���k�5Qͅ���n��:�M�s�_u�8n���+�i9�ޅ)������(~{a|j��?|KT���\^\�%tz6�҇����3�o���`�\s�����ۭ[���>����u��f�-�#Y}(����=/�lveE��S�D��b|�t8uv�
z�d�Bx�4%��^�+ݠ�d�\F��-����CJ����lyj} �Jڧ'j���*�^�SM ��^��%�[�q�"MJG�E5��{^��� W����O���#�vT�a�؀��IY�?X#'�nD��Q^�� �e��S�]Ma��xȞ�n�*��Rz��R�h �AS��QbQ1 �W����m�@ZLP�
N�����-ޜ�^ͭ���Oq�FC�ӵ�Ɵ�J�;!����	v��v�\!��G�`�[п'%��pP�%xX�"��}��I�LS�"N�C�۩4oN������-1�$��RY�:.ʴE�q�B��R����5��2a�&Cӊ�fgZD�g�6�oʼMi0
ka���7֔���9?����C��e���e�>� �)�#d0�h�:E��;�	��J�[���[�F�p�΃0�9�!-Z��٘��)�x*��hҼd<��e:�d���9w�����y͆����|BNn�SޙqZY�kWc��t��L��Z�
�M���/m�	(&2!�'�<x�$�F�a��cӧC�ȱ�M��)< �.E�;���+���w��A!qI){���Ff9��G�"�(���v���oj��>L"%��J���v)u��C{�4 �~>6��ر�Y����#%��ėoB��&��BE����t��=�3�ir���� g��Ш\Ku�G0�J1�ۺ������҅h�}�����\�����4j�T��x}QС�b-Ap̎�����5�)�-SI+l���S�˻�0����V�S�ۃ�!��O�c�n���-lV����Xm���gj�a��Rʧ����ua%���r\�<�Z�{ �X�#�l
�U� ����Ƞ��栣٨�[\���/�3w#'0ꐻ:��W�C�q�@md�Q�<C�Ƶ$N^��Q�PwDz+���3�Qw�O�6D���gtG���ak��G�i+�����]���,�ysl�l:�>Um0�	�X�	��ɟ+���E~I7���'E�u6՘th���]�+-A_�ג�Ueu���Qcг.�H��fq����&��� Y;a�D���ٱ;,������*����zw�kEZ � �6��3%cn�W�?6��P��>;9_gx�*��"�םZ�H�U)�DB����v=Es���)���hel�H��/zw���y$��q`���@|�Ľ�>����nR�W��i�Sp���NN�x��AN`N�����*j������ʤ����& 8W\�Z�����*\[�Yo;M��n�����5#��ϓ��	Y{>��X���Bށ�r��LVM�q��0&�k�2�~95<vA��H�t�-����j��d��:˫PD$X�M���(�����T� ���!c���}���R��9$����mb_���'3j�ܼ�oB��
C}��gy�����\���׹��N��I���l��)��VN�Αg�UN�����_pCxS�j�T_P<n����1�m�X�?�q��\��`I�O�}��Sl���D�:�u��;�lq�3�M}��;ft/���ǡ1��~ ����5�A[���7 ���$YB�����^G�V����ѯ|{$����*�h�1���-z�}|=|�x��ң�kv0�4��|H�_�{-	¨@�{��}0%�D����:�,�����C�r����b>kCSB����-c�G+V�m���Q 8⪵�,  5}%��=GE���i�Oj�'���^&*�_B:^e�x	lmG/0��FA�0�RF�l�H�����'��G�':����.�!ъ��~w.9sGvq�s�'�Z9E�𒱸��=BN���v���P�'\�X��H��S+[Z=�Þ��"�GV��00$m��E-�<>�H������9��\# �[(y�x�P"��p[�E[��J� 2����B�=_Fy�F�s�fޘ��!�ӽ��4����^�ls)S��h����C)�eǅ�of=�;�A/-��-��'��b2i+sI1�PĒ�b\���:�A\q2T�~�p �W���_�ͯV4�yrl��f\#�� ܘE���9&�/)fI��0�vi:-~�Ǯŭ�r���_q�*ҜS�7�[k]s���S ��y#��;T�B�J@�S����#�nT)!9@7t������� �T�=�s{sh��������]SJox����{ցΉ��-A<r�ސ�{�$�T���@��A�e��?�ܾ�sA����2�x]k�*�kr�����c�7���%h0ýP�L�%L�/�$6�B�MŌ��^��k�=]nt��ݮ����9��)z���s��8=�����ci>m⛞��>���V]#��N�f�S�cdg{|WݖQ���^��1e����3������>]	Z�A,�*���o�CyƿՂ�Q�`���E�ߞ5�X?�w��pЋ⚔����1�Z�1�3���c�!L����0��%�Tg��.$7噑3����En�:t�2��pt�C��M}�r�`�bf�g������<B�z��*!h0�=�B��R�g�%h��ߧ�QA����>jܔO�>�[9�{�M<?�j�[���S5I�$R�g��jk��~{=QfVJP�*�;�^�9�맘�a]�G����WN�i����w?�s���-/��*��~���C=��	 Ck�����'@	��oij��JW`���Kv�dD�0��*x��\��/y�v��7R�u-F���2a�9K�n��9�n\���(�rə���S±��3�-~��a{��I���zw��yWS.�P���Ub�{P��v���ղ
b����(�H�n��R���z��F�7��MҋJ=�gG;SZ+���!��$,g��A�]�V�ջW6�9�V�hW�y
�ux~/V���A�)���_�X;j��M��&�@_�`���� 6��>q�>��6n�&I~���eg�Ⱦl� 1��2ya}lt'R�Y�B�"�W�(����S|Ƣ���&+J��)w����`qBo	�u.�n[�&�Ef�,�L�i�4�>+ߐ��
����uB��Ӗ3���o������L%E�?|�J�����IԈ�DycL���瀅�י��g2�a��H���|@n����c���뜱��ӕ��[Sn,�E-��.�E������SL>|q��UU�}ȟd�5D-��eҮ`��*h����Kq`�Ѥx���R.T�"���B�#�I��
�jV����n�?&9U��9%3a�ֿ�F#�*�3˹T�`�@ �s{=^>��)�Y��O�.�6�g,I���ɰ��eOS�x8��S]�3��4�9W:�_I�^����'�1� ��s�*���EK��<�m'�R,��-�yhr�N/+��R��_x �e�����͛Om����a�;�U�Xv?v��j���a����a�a9@`\%��Vbb��T]~\Cۭސ
�;�f+�Mn?���C�E��a���(�����i?�u\w����knc��ؕ2������%Y�۳��Y2�0}���Q&��
�˙�ǳ�`쇂$z���JLD�ķJ�6�l*���XO1�܆a�u�K~F���t�@ZV
�[ִ�L K�j��@�:�/ ��-�b�5Tܜ֢+��4M��D~q~�z߳�������>6"��,�݌^�ێ��,T�:�
��"��ۑ6G�4l,����iyA]%uܖ�c��h"ҳLqVƨ�9���b��}�$>��>�E�=���'X�-'��x�:�~t�SsQ� �Pnou��d�!��ҳ:�g�	џ�����Z�:�p¦�!RN�G�?�Q�͘.�U�#zWwmxj��(�a2r����׌��\�$ ��WQn�C@��E�ك� ���gͰ�7@���q�m�R��w:.���V����*9s��fP�c&�ǲ�N<Ś���@(f�Z+�)���gB@7��e�����Kp�u%s�rj�]�etɨ�=�h��|/s��6�Nd��o�x&ߊ1�����dME���[}��^��P�* ���=����J���� \8�=��($W;��P�i��lA�I͊3̫t@8�+�a��XF)J��S;a�b�+>�0˞���П��{`�=��,�@1N%H7V���pV�~gX
B�!�j�V�>�#���f�Nr�.�{q�^;����(���c:��-X_�6x�P���֠H��J���?�y�+~��AN�
�*�'ټ�	^��5Ź&�zI�yp�V�"�}x��T�i�I.�nbC�R���A������Z+��ue�����s7�~��uS�[]����_��S/�c�Q۾�e�bC�i����I�!��s����^�k4�@!�h�P��Cre%(3R��A�m�m'\�M���0&����&@��QҍE�4�;�A�O�O8
��1�Y����c�&B9v�P��h�2������ۄiRk�4��mu<|�ј��#D=s�J8��3jO��-��w��B���j�:
������s�*z��ō���k�r'v?�֡��lR��4��a#W*1�t�OM��W�QA>sk�/�Y�'�e�!+�cu̥��w���*��Rχ�;.�6"�)3��Su֑g��L�giQ�!<=� OX�����f>���A,��]8��N�^��zw	o��r�IΌ�=%�IB�̬�RJ#�8-�T׽������L�se":���r�ҏE�ƪKA	GƾD"�L�v�d�ʙs���i^��"�����0ܴ촭L.4$��<:g��ˮ��	@�ԥz�Z[~��b&��b:���;#���ޠI�%YLϚ����EI�����-f��l�X�z�F�'� {x̊�Nk�ZY��6W8sܣ\�����Х_�L����Z�~^���C��ͅ��$־[����R��,2��e�Ή�������	{�}'P;��Aʝ.�0�SIQX�6���1K'趩�/af_BX�![E�T+ƌ��d�?�k�(��Ȥ)�4��c%�;�Kx��:)PE˃��4	9`���qy���;�}�h�����y�)�>�y��	1��'��Nk���K��(�v!��:{�lE���Ƶ������{>9�������Ǯ
/�ʠ��s����X��ZL�ܪ�L����G����(`s��r���,}�m��%f�q�/c\u��ai�ϗ�JaD�t�wv׏G�J��,��� �$�

m9O��C<������IR!g�߰��dT�cI�&4c!T%�zC��'s�j�,P
ת1��ؚ׵vc�Җ�[�����f��5rsA�x� ����Q<�6òcL�l����5�L��]�G�@Lu8�r�u��:ںi�3�E�V��y��o����D@/�O��M�g�'�Ls{\�PH��k�i�3d��J<-r m����Hʞ��Ը�\�_#�Q#@�㏙���(C�P�;W�LF� c���J����&���Y�:�m�y��u��v%vgms�c��oT�C�$��$|Uw��T���.'�ݚ���N'�3�A�K�����.�hZz	�0�&߀���8Y����	r��[/	�Č���I\+�W�w���y��D���ΰ5�����e�e9מt��8�O�������X�U��?��N�lW�;�ʚ0�2�e�
�����q���W�$h5���;�!m�Vd�2�˜A�B�-��VZpv�I�Ѩ���\�����a�}S��V�v�˼\�nl�\����{`�]���7Os�QbLt�3/JB�èz�X����â�i�d�.?�0Jr�ˈ�\�6h���\�JQ�uQx��[�t��&�\���}!+��"[2Fxc�;7t���u��ع��r+�oW`ߢ2�m|:B��8�JF���W�{��,�7J[�|t$B�O]|�n���R�8-�¶y������y�-g'PLA��sU�4Z.������r�E����h�����zV��3t6 Nd���x�~=��t���ЩH`VQ���q8�O(�z�U�ʃǈ����ʴ[JWF�y�h޻71l�{����T
�Akޔ>{:���;�n��3������۩#,��k0�%�� ��&���pn�)7м��y+��6���K|��U�JU���M��R��or���9'H��{!�����/r����$@L�q<,�vsx	�iϼ�~��k� ��3	�Pj	�:@V%�טj���  `����*um���I�-��w��fC�����)t|P�l��f�$�xe���w�����d'T~i��k�]gsD�wT�`ȝ2��Uɼ�n�>��Ņ��q#�ۈ���]��!�8������~��Bs�;�*&�4��3W�k`&��k�5sޫ�i��j�M�/c�N�Ya�o�ąм!��?�Aو�#�왳|΍P�l��!��El���� �2I�1�P���`v9�wA����}̈́���}۰��nRɶ��^����FO�n��7�6�1�����c&qn7��p�_�*�t�a��_heX�E��*)�X��c>H#�yH��Ͻ�Ka	�ޛW�w�I�j�� F03��Ǧ��HQ,9��Rv|���`�ҁ,�/wv3�5��p)R���iuN�^k�^��@;��2�>�.�.��A2��m�m����1,��%�gqjQ�P�^�U�QGU��S�0`'�E��,2�l!_��~c��{����ꉒ`R���7���W�+�(�O��wJ2YX	��!tN-9���ς�����7���ϡsrȎ[��m!���_xdX���g>YU���������K���W�]��l�>���j*׷���23F�#�8Ӝ��cZ���ߚ�nӋ��JM�n�9���~WTK8��a:��5�ċY��!�[^�^�v�ޔ*M:���4��dR�'�{/�M��f�'^�j�	@I�A�ߌ�Jā� ��5�u�;ew��񯳽YA��Zi-�~�٦��&���~]=�}X��d�hr]�Hb����<�H�xZ�C��������hz�m���I��vZ�Q�w�כJM/�C�:����N1#����|� )x{�'\\ CS�#*FU���~G$MB`d������O$���@�#�]d�f���Ү�=�$�>|yV������9b>�w{��b�m���D=
���@#"�&'��A� �9}͙�J�.��/Lk�,��W`��LWʧ6[�pJqt�^�1)��)��m���OM�=��]\>^E�AHE�ܯeB|�����92�GyH5�߶nb����)����G��i��/Ƞq��׎�c��B/��:Lh����=Ms�#5����w7c��&W��9��c�������ø��(�� f�4�:��pȃN��(X��1��MY{�ph0�ȏ��c��SYO{ĝ�K���g뷢���3ң�S���4�ei<�f�I�����G�A솫:Z!��� و�r� @��%�h&���\̜��z�6�܉��`ʏ���"L�l	]��_|T�a��c�L����d�3* ��/S�7��s�z�U�[��n���}�P���OHݘ�z��1��y���\�) 4��E�DX�K��e��}�#:��V�m�X7�5I�e�����k6���Jz��p)�¹�/0�ҫI��e���_b2e����1e��˙���xw�'�D�f�����!�H.<�n^3�
R^%<C$)�� S�2�j�t! F&�����0g�e@q쑖쩙�����'��3�+�ů������ia�N�� MP�M7(��?�-�3L�-I3G�H��N	�.ڇ_�:I��;N���H(�s=Ō��˜E[�'u��hL�O##���)�$G�k�-6_<�Q�P����a�zNR����&�3�N�4*�4��6	���럓�Tt�Rs�4t/��5���g���O��fa��2cT�aGE�V9�k�8���3cn}��+�x��c*��/�e��$��G#;���*���.��/���;w,+�����q� ���w-*^�b2��k�˂�N1��8^��p��h��F��l�)���� d�>��w$��;�<Α0�3���^�N���Ԕ�=ó�0��5�?$e�"�x}`D#�@���r$��1H��5����$�m�%�+��_�R�ʳ�4�Z\\������t�a��H7��-����<�[�v�����i��<�`<bz6D�	�Wo�o��q�~��z��
7"J��vZ>nB�ņ*�Hy=�7:L���,�U
����Dwa�������q��߽����Iv�Wq�����������D���̩E���wF��^�/`�A�*���C٩��^�7۳^-����{�{�zr����*<��!*���HDЩqȫw��t��nO�����j@4�r?�M%����1��Ke�d�������m�e����`�"h-p����V�ro��~8k��$�T���x�k:�ّ�2b���NI�1��C#~��\�z�Ǯ2f�k^o����'����k�ɳ���ob���Qb�*/����G��f��A/'�W��+�UN�p�!��-� �M�sZ�N���>1[�k��ڃ��h�vj8�վ����Ϙs#��������F�u�l�X��N�b�<p�F~��5���Z�lY�e���v�/�>赴|P���wd�d����w����X�$�ϐ��]��J�ʲ��QB���	a�a�Li9�f��?�[x�s ]���ퟭ/�pPަ��%�v��2���-7�p&s&<sQ7�Yq��h��X��uI�������N*ܐ�N,��S��kY����*��%G?��xxn(���L"�GLܡ�B��I�-��W��E�Z�6f��߭b��H�֚��4��a!�����#]�Y:�^���N���*��'G-�Bm���M���W����:��3R�W�Q[��$Wb��vLF"�I.P�4�k#��?�,ݜ���}ޔ�o�:#����ԅ����3��Pp��,��e��^�>��~�|7A�l��=�ϟV��N������e�ﵤ�X�:�G�lg׾*��_���i�9��!��] B��e4P�BأpO$�>V���p��bŭD���n7~3�_[�Vf��"��b���R�d	a��h�^Z�VǷ(�?�����)�7�Hp=�=��qEu{�2���;�󆸚��&P7��K����kn/��;����_��ۧ���ĳm)xl"E���r��B:$	}Y�*~��yZ��XCjp��e֊���	Z��/��e��C3à#�=���xW��j�BNH� v���2��)���B����z�1�E���p�B�j�l�}��+���	�����w�%��>�%������a3����l�<�QWUP
�$���vXz� gq�<c�Gc凬�K������FR�5É��dn*�8������	/j1��hn���*�E�?�^��0�ͥ�/o�ܯ�O�1�����S0�F#�^Ůٯ����O���膒)���ȸ3OW*~�۾����v	0ꀧ?t�R�^��"�u|��R��V��U�<�A:��������t,ٓMB��/u����	M[�=���.}���]O�2n�dT�;�:4a��0����P �8�$�k���Ǝym��&��x�Ӓ����E�i����
��& ����ӼݼZr.���<Jߧ�`����/v��)�����388�G1]0s�^��T&9�<\2���rx�-��Rq�<A�$�J'��y�?��2k-�B�=,Mp���E{�R��c΋����$�.����Z���}1���[�,\"D1-����-�P_!&��=�P�	��@W<4����>30Ѐ�o��o�%��y��:�u<Q��?WfJMTjߝ�>��^l�E��"��["`}=����)���h��?)x\:+BZ5�j���>�y��sl1��~o,�(�uT���~�VҵI<	��ni'�z�����mM9�?�ďpTQ�
�wf�N�~�%�r7�因�I�e��3x��h�B�2�G&��5�F��{^to�Z��&�]����b����m2kR�"nW��P�Ls�s��SC�:Q_�Rڟ�D�#]�� N��o71����^u�s�rN�S�EȄȡ�hq�%����No)��#c�� �����D�:)R�0y�)��n��v�ģ�QIX/��ْ�Y��RsY�Wk:�#Ň����q�������u8���]�Dj��C,���c�oe�yGŁ��̳fX�@"	�K{ϸ����'ѩ�n�C�C�t�(���=~�Q�U��{aI��([�� ��*�=�[�5b���]���
���%��04ph&��G��^�{�|O�'���]��q8�������E����z��_���MdV)V/�-�o"jh�iF�����X�V���G|�Z֟�H�9wa�e�R��6��3���eay^7d8A��8�,Np����CT��:��~U�x��fOv">9�5D����-����=�Qfg��JC2�<�o�WS�L�<�]�~��Ev݋��M+���\�3�Αȓ�+LD2�=I_Ud-WL'壟(��QhU4��&��N���U�ǼŪ�9��ؔmL�d�/v
�ξ!�ǆ���$S��v^�T���*B:�6�> ������7E]6A�'�j�23L(R�i�T���˴:�-�$�sD�'j��[X���#B17n����+�n��sK�����|��^��|��k���"Ǐ�U��FQK��?2%IR������2���޼#r���IgΐNdzd�֎���o@���4#-aK�?EZ�GW?\�_u(tָ��K��2�8�d�X�V "<D0��o�G�MuOT��=<�a�*�UJ��� ���3C0�y_��.N�奮��p�|��ʐ��nfV��~q�Z,S�iz8��.�EJ�x�n��{���]�� 8x֭ʍ����W��2�/�hep\�L��Ca;m�>��ڼ�C�T��j9�DM8��-�ǊaWe����T*Yv��7s�*~$�����>�a�e��A�����#��P���50�7�p��(w\��W�dȲ���8�E��[T���+�!�A��8�cu�ӬX0��;	��3���D�*,�݅}�X�{a���H��W�|�ܚ9����<�F;�Y��y�5�Y�T�ҳ)Wi�B>�l~�$������ ߆#t���kg�����hAK�Zv8��k�L
K`�F��2��4E�jx#�1:(n�^^d���٢P�cr� 1-o�B�R��BdI{��:�N��~D�5�l��X)O���J��=�86��lU�@5�� �������Rْ���ez��g�٨/̩#�OR�:��i� `�vѣ��5d��iGNrD�6@U����A����!H,P�K��dI���1;/��8�� z1)�wd�B�����kR�`ŋ͠���!|��<������ �_o�4D��t�hky0�X���!����j$'������t�>ա�*,O�"�.��#�Acji{g�d����a���%mC�_pc��17���"_���O�0�U�p� �ePt�1�&�WЙx�7���%y�+Z̓۫�Ӄw�X'�~�ϻ�p������[�T�WO��8]�5���#��ᮄ���0�kCu�Z&�±h�և�=7�}�����d<�������8ᧄ��Ϋ��)��E��%�^�� ���k�+8�{zB���G�u8�]�K/�:�J0���V%���k�x�w"��>�@�|�Xj�I���	��(�Lnj*D��E�_�*y-���͎�, �[������GK���>��s���s=��0e1!bόz�r���t�q&�:�0���$;p����$".?��'�c�h3y�Ae�>_�iP��.�O.V�Y���"����ڤ���"�Ҡe�fR�Q!N�B.>�J{7	�^�a}�yJKN��ޤ�F�؂W�4��%�@z�`Ǝ�9QFAB˄�88O�/|���<��=b���J1�VYG�})v~t%\�[�iR`|9wo�v��nU��1aq�g�T	əT�8��߳@��;�M?�G����0�䆪\R��E��UO��2��u��l��S�M�PGH�_倱���7A;� ��СvgX�w=��$��X�f}c��1���E�>�z�iN$!��=?�!߄:h��d kO��ƭ]���5�r�j@#�0i�1�l�����A�#�!��.��p�̓(9����<hٳ�v�R��.�?�z����2���M�@M��V����J2�b��`�	Ǟj��ńɶE6��y U%�^01]I�F����;}��{٩���D��T����u��`�I��OD�k;���3�q�V�������%6J�7�D��,�&f<�[�X�'4����(M[k%ڀ�[���1���N�D����>�":4��r�R��M�&|2.��<Ep�Y���Bŉ��T�ޝYXw��qS]?��Hv��<g(��ȎĜ�8uNjQJ��?vOZ�=�v���xg��`�!�O�#Q���0I�ʱL���h���{y�)�7ζ�Ū�]�g�-k��I�:LKfS��t9���v�9R4�{��;��>&���-kO���E7�s^�F�5�����,�v^=l�����a��yS�ꍾ�a��{|�hR/kN����L����FSwdu��,g�.i����1�D���¢�8B!��W��ֶsZ�_��a?�Moa�+o].���C� a��{t|�~����G���u�^Hrd�b���@�����ڣ�贇dYq�Z=
8ί�7�' �	Dd�Єu�U��e- ��N���MV�0�%,��V֢�IDPV'�KKq�oE�.�'����I
\Q�D0%�=a/�#�!|R����fBL��ܙ]�z��b_'������o�'�зK�\0 {Ls�N����`z�Z���$���Ni!��]ͤݵ#øq�V�0U	Z�,��7zu���
�L?�ķڿ�L�c�I�x`G6p��B��c���0��t+�}��Q��]���L�Ҕo��k�E�{L$g�$���.eGo��G��v�NZ�JV_"ό�2e�IT�]�4!��[��l7���g� 4��sRS��oP��v�*����s>�n��	Ufz���d�E �4�j C��-C"r�ar}H�'�W�J��I�%𧳆��Ώr26�:���:Y]��M�/����$������ަF��R��(Pt�-��4- ��C��I�Mn�u%3�{�!@T� �z��kp�b��"���o�O�$�dI��)�=�·�
 f~�y��y_�2�h5�\�������HS���PD~sJ:`��6�}��b�d@�<R�xMR�o�;1!iy��8K7T�<�班�7�y	$�QE��q�J�g��!��ǫ4��o��4�	�P�����[W�U*��,P���?%�Ww>�E��US�����`� t:��E����A�x�z�n����IҚo��mrߍ�Ϊ��}���D�m`������S3%w��W�okGB�P���|����У��	�JR���y$�;��H_ ����~��2�AN(*��pqʂ�1#���C^?���[��)d�������M��6�h�r��e���MI�$m�/Cį�a�߂��jYXa�3Wd����W�􂜧x:�18�����ԕ�4��&��U�\T�'��{�\���k��+ =�&��j�Y�76�q�g�񇆅��ڑ��'k�|-�.���
�98X��|o��I�1�
4���#'_X�V�z�R�Ǒ�H������7��JiE#������W��<jK"�u�fY��%�^q0��H��6Iܦ/��}��f�"Y%�$�j� -�!�8����b1��7�nߚ?�A?��F��u�L���&u�C�,ʘ��f��8,B0��n0�dE�^�ſ�Ń�od�����=� �_�j�����4U$W���!��e��eӅTɻ����Έ�Sg@ri�wMB���K��7��"�4�]���Y�	4��<�]k�vG����1�D��"�u�s�]�|��4g~j�:����|̈́D�i��ZP�&/�?��`�MS0X(8 Y���֝�1��G�,\Kzu%�d�E�C�j�5W|V"P��0z�㽿�t�{\���</yL�,�"rm��zx�����C؜B}z��-=U,TG�{�)���_�2��*��Ÿm	�L��7c�3��4+O��c r�C�����g���y�y����$�T�$3��Ety[v��:���c�Rx7�p�Z.���C��H��Sb<7(~E:���+����:�;j*)�t���O&-�Gv���[J8��"�J�ym��dp�,(|�N\�>���MV���
^r�E���`��r�q���1�\�: ���־]�F��
.<�����KM��j���?�3q:�5h��l=ngo�:��S�T��yJ�[*����D��]>��Q��T��\�<���F�_]�H�Z���z�c��x$�
2Eut��΃~Q�-���+��}TBz1�#���R�M-yH>x���:������k����վ�~���\g�~Q.��-�D�����F132���پ��/P|ӯRҜ'h������,�Rpߝ�k�Q-��
�4Gn:��]�����b�Sw�蝴��s� ��#�XbF���<�?��vqV���v���N�z/I����E�Oڮ�3{�V�m�bj�����ccK>���?T �Ij��r,[t;�^	vv1'&�gܕXJ�e��-�-��n�:aD�;޴�0=�"Ζ�;��
��P�����7;i���p�ÿ��a>�KI4~v�n>��Ӕ��L�����)��T�!3�?�^B��Y>N����cH"	��K�m-�<�#�����/T��_}���q�!�V.��ZD�u�JpulNA�/��d�����s�YxQM(��q+g��i?�j*����Y�J+K�ʜH* �qh�g	�30@?� :�-��C4�[�l�M5��2Q�&En��P�8��W8��t�6�{�s��geT���DۂeW,���:��|�hL��'$ؘZ����[�>�7�=͂���(p�n�P�i��t��܀]<�p̊
k�0�x����ݸ�֋�$y�	����?��g�&?�i��
��R��0��3��Q��9}��5�i�[j	0���K�8D����B��a��fum�\�)��D�U�X�7Jg�#�7[�+��4��!e�,6!ƾ�	�o�X
�CL+x)�x����DJ�0 �����9L����-B��U��E�YL5��-��Fv#�A�+�g�8h������W�("�+^Y�9���v�ס�M����� �U� ՛}��^K��>���:�/Um�-�z̸%$t��Xi?	I�ρ!�W]�$���Sj�<�71��3U�_w�`tpi���Ȃ���m-�|�� #���B����r����M�ˮ&Ȝ��T�'�hd���7�`�*HfGo����tMYg�D#��4GT\�D���7.�$aV{�r�C ^�����~ֵ%a��v���ZfH�O������N�c�8���!�w��hZ�\g e�H�L�x�R|��m�q�k"����0���.��@�`�|i;��=R��\C�8�$��.ӓ4�=w����D�����C��^���־VU w?;E��<A�"Ye^��Gefv�b�q���te�"�e�R"�s���F�Q�����85M�Fhm��o���G�ᣫ�B�JW`o�I�Vl�	���A]d5�lX��P�u��Y(����	�=~�a4�I���*�Ȫ��b�o�V���&�]�TT���+��j�B��}�¿��횮'Ipk1^�Z�b��o�V��e��w���� �RV�Y��W�#��c.:Y����Z`���-�3��uE� �
\n��' ��rhEPo�N�Xݏ-?�(��
lx?*#r����qƬjt8��(���G�`�dRR|s��A�]��¿WI/U$zֱ�u3&f��Zq��↩%,z!F�$�	�f���,&m��Ս�G~�[�Y�ա���;u���)��G�{b�3��ҋqx���w�l���sx��xh�e6�%��-���
%z�u��Hd�X݇��׆ �'�ҍ����
D�����h|�����!JI<� y����4��y�F��-�����A^��UzS'g�љ�0G�w�%�k�:m�s�H,v�[�YE�����hI�0�����Օ=�$j-�%F���*�ѓ�
@z/�a*|��n,sdiQ�uE�s� F�(�~�.���[�ʔ��t!<A�H_~/������Ƀ�z����jW$�&[@GH�s��O�z��)!�:��SS��?���y��:�{�,���rI/�ʪ" 'ļU����cG[0C�=��=�W�d=*l�C7�$;F�T��5�1�t���H) �)�ї)�2M�M�eڃ\	ztS�C�4�D�~�+��P���;�
���X͗�MSZ�`�Im�[���(.*�;0���J}�={H��֐u�/83��҃��נ?��%����'i$m5*D��0C�������v胲�k�����,ͅ�3i]�����!P�_N�u�8�|�)�D�v�fe��ݛ�5=�"1�X�(��I�/I���}���^��9�ْ�z���oxO��h��1�9��ρ��o�}tE��?��� n-:�99��~��zl��Gl8Z'죖k�$8�fW�Dj����[}��ы��i�4v��������i��n����a���I��B�eJ'��Cg�'":��t�%G��HqQ�5�Z5��vZ�׭H"��gT�\O
���T$�m.w$"EWV�m�G� �Gl��-~z�r蹲X�������/~��Z~H^�o<�_l����A���TA���*�K�m�N2�O���J���c��.���Uw�Z�E�0fL�:NT�X��ϼӠ7�-V��L)�s����V�!��]�9���J��Ml��@�)����G��Jr���#p��oq+�tK2mmTF�IN�&�a�(���߽��n�˘v靈�/�t��,3��!�<;���X�!�XKd��/'�&���$�n��_?u����Tbk=��&(���ż-��/�}[sGr�]Pg�R�Х�9��R�����=���+\��zBa���g��ohD_O*!��q��4=r�!Cz-T�Utq���e��P7d�O1��F7'IݞC��Ej%���-h�)iܫC"�ľ�yɮ����ͺ��RPq�S����S\)�w{�ڑ!�B�*\�Nr��V� R��辱��G>&/�	c�h��ד�`r68�%z'ҿQ@%�p��cLs�qF�k�3U5u��S!g=�w�5��u��B+"I��Bnh�K㶱I�2�:���J֗��-N�5Y��m-��<lD!Q�cM�R�"vt64���M�=ɩ�񶯊�<�s�:̹���/a]cBɠj7��9���w�ԔS�>3����O)���|{/*���=�9�u0+��'��'��sb�ǁpB#��+	d/�K�0N���.�A�5ы��;9�+��'n�x�?��
�21⛷i����ۓj�;s>�wi}8�^xi����m�HZXx�H���L�@�ݟ����h*=�� 1�ܰ-�����܅,:t/d6��+nP�5�(5i:JZS[}���юhIm��.6
#^���T交��$�6����K�<]?0�s�;&b�?�����L�[��������cv�.�3���r��ET~�zZ�������{���2AOXm��!��۰vB@���!�jjO��w,�:Q+�Y���Nh~`��I�N�����r���!��Na&��)t����0����{<�Ө�(@�$���F\�u�V��0��u(v�s�	�f8\��Xiο�55���Q�}�Pz �EG����D�m�l��D5��6`�o��E4�� ��3Y�3���u�9�cώ�7���u>�=�ű��w��P]�tk�E-y�elU�5�%-yUv|�n��\V���Nr��e�2��?-4�=B���ޒ���Y��6�k�Qw�l�G��
s���Ԩ�c����xr"�>�G�(9oA��.6vz�J,kj��s[j���J#_Y̾�
K91^��j��@|aPbR�IZDV�k���i#���g���in����-g}�d��5��h3��e_�AhC��^�q�%R�������.�1'���>ū�#M,�����z��L{���5�ä;G4"v;r,�����B
�V�oŨ4��|,]����$��lE��0�'�{�xs:B�
+����|w?�]o���2��m�����^I\�a_�K��2��#(�v����w(ʁ/���Wr�[��Vˈ. ci{�%�~H&���j�9J$�X���؛a.U!9�!|�˛�&�'n���뾒.���z���+�_�xJ>�?d�!"�yj)�x������������l������03�E�ˇ���C��lxڴ����F+��dzt�q�!�����������L��^�3wteJ�܊��P�ü5S`w���=~CRq���o�+�Y�������.�Kke
�\������z en-��~�G��9�߹�,Cm��m?&Pڏt�̍B(��c#O8x�:a��4H.��N��  �3e/�ۜ�} ">�Z;�B�������7��m�00�ۛ*����w�hي:0JR��C�eY��P/�V�Ht�jm�X�F�<�/�g(߼��ʠ�E}z��k�7�Z~�8�Y֣0gߗ���F?E�/pڒ0�c���C���*��.�bo�sm����
�o�&�]�y���t�e�1ޓD?,�$����GxC;y�"�!@�����猫�!o{9%b�5�x�栂�� s)�{���)�X!J����=���ȡ�rX�	�Kuq}w�w[����Յ9B م�z�ԗu������#r���*���������#;?�]�:��(�������*0>��k�5	b�U#*���6�8�WĄ��{�i�������jC��ḁ�׮dʻ|A� s� [_u^YE���d�^�����n:��l��-���BC	׫P�7��e��Z��}�������v֒uߌ%_F�5�Sњ����*���ǜ�����E���1>מ�q|����Q��1\�u�S���&а�G9�h����7g���T2��#R���"�gB:���!���J�nu��v�%E�0�},!-��6�`�U7��{���N|b	�9�"���}�~)���ƍ��nO�]:�檃��GA�?�9u��s��B�֡a";��B�d�~��M�ַ�w���c�#76˼������썓�������wJ���2
�?d�S����S�B>m�@�W���QA���{�&sF�ַpҙhO�������2,&�5Y�lO�$����bb��>Y�$n� �B�����E"�N�C���J�ΕFxPBڱ�\� ����6�	�h��vwU�h��`"�h#6!�}���c��q�.R_��d�r����}֎M/�{���E�Q\yD�� 9V&u%#j���RN_�|u?�[��p�z�p0�C�z5���-4ū��T,|=�:���C�o6�.�ʖ8�&KU���ˡm����U@!e���i�(�O��� �j��h]  ��L�Ze6Z�K�B�RE8�{�\I�-]uPДp8z��xH��A]@�m%+1╚�s�d&�u����i�����l�����\�<��yO�=�#�|��`�' #�)bT���X�)�!����v��^�ΘZ���	կ�k�O3d\�f�`9��d1����,��C���4�p�ll��]���|
|y��Z�,ay+�ʼ0�z���i�E3t&
U|���?j�+�\G�������ҡ�B�?#�����la3�Z�d�T���<W=�9u�<$@V9�f MrB&���R�齷�rV q�YWܨ��e�wJt,vHo�6k���ZG�F��y ���Il{v���v�6m����4���B��Ѓ[�7�D�/��J����W�ľ�9��?�/|���u�\�Jy����D�f(�tG�����7�G��e�"}��/�Oޏ2r�`9j����cJ��I�"@��ң�o�j�,{9��ܣ��'$~{v�Й(����) �����{f��9�m�%ػp�jo�܂y<��Wv������C�"g�S�{▃�N]b-�ǝ�1^�6�S��>��F|Z�АZ��-��8v*�����ס����.�#e�t@�ei��g;p�]��/�^��u��x =V��A�sz�伩-�{��F���4�f��&�3^��hݨ�@�+�nZW(����@xl/Q���W�!'�X�bjI�u�d���w!�l|�1}�yj�����[8��~X`sHSe}��ʙ�@j���"�i���6���\H�o�⛖LߏQS���ZF^����}rugf�U��p��Xyo�pWI���myR7u{���I[%�{���]��z@`������㧀�q��,�Vq�����6l*V$���������Yr��?�SAV��`/��@ؖ�.�g,�����K�5�ԌN?K�A��>W5|8�o�r�haE�R3��Ъ�Ts/�mY����cѥ�u��pf>E�,S��_J���,��0�����jTiR�v�������1hf�fE�=����)��M-f�e;�q�X� �<̥�UY���	�)`�p�t�h�!�rx�Vj���1m�%G��0����l(| O������wp�-��~����];�T7���f}���ޛ	���JnE\('��r�DX��$�䣼JT�b�w�E�5Tb;����5Ԛ����z:8K@&@]X�X��Y�.�����Aٱ �amp�!aȕzUP|~+)���ʃs�����q)�"�*�r���oż�N�� -���b�����mh$�Q\�Tu��j���GP��p'�TQ���q�������p�i+6�O�w���������٘R�D�`�l�]�9��'��-[/�B��L�-�~z�{�[+���E��$,�	Uȁ!jת�,.�Ѭ��5��B1�0Oa�vӸ~v�[���3RR@������Qz����X)��J�>�$��.���Y���ؼ9rG�MrSJ�f�}����2|vF�z��3K�f: ��?�<�|D/�% d�C97\��sgbk�K�{E��R�5���3�ڶ���v	���ǸCy[���G̱[a�4�߂���}huu�Dh��~Q�n����|F8�t��B"�� P���ˑD�be�cjP/�f�@?�z������k���	G�(��y{�K�2������X���6cb��ɿѮt�~�nm��ŵz��K�>��Y`��R�6�+{���_S��1E�rV��V�#��%�������%�=�\h"��wpV��y��3�&V��Q��쿌Ֆ[�bxWPHQk�Hz�$ $Б��;̀�Rl�MB��4fxҫ���)|Q(�Y���ctm������7���	9(��ȁQ}(��c�`���v�U��[_	ө��`\��v�� �濣v���m_������;M%ȵ ~0�B{z�$������)�+���9e�P&s�E^�P�pP"�"4�L/Z867v�{��ظ���2�0��ΫK�}^x����H�	u�4��Y%�������(�UL�w�x6�����1�8���O`��5Ksn���c�9��K�K`�d^n�iב�Y8�^�ܳ�S>�M|)0?�\f���y��3.���-m_I`m���`dO��Z!��ğg���i����ҥ���8/`�z$��Q��Fd�c6�Xp��<@��VϝZ^�ՀAZ��%6��h9���&@� ��Y��!�������R23���CJ�v�l�%IB��c>@�$ŚK�(]�d��9��Q����{l���?�$ӊ�6�H�1��ق����ђ(;���h�q=a��AQ�\�y�/�#�Ο=F_��rƘ�����3�;���D�A��y59�'��-Ǖ,�����������0P�1�YXp]�&�߮�,f��A�+�m'�?�4=`��Po�mMu!)/i�蹉ƈ5O�O�8��Qp��� �X��/��b��&�f$È��-��o�� }�P���q�W]���w�^�=��Y���x�[��5�N��{�%�����*Yĥ����\��)�{�&�b����5����tf	ʷM��e&�c�Xu��7p]�?���-���₤�~|4�Xv�姀"��2�.�N54����o�Ä�805Y��UB-c�j3�]`%�/�y�7aޣ��,t��������)�(�Zk�9TZ��I�s��"�F�����7k���#�������߅�}���{�w�n��l�1l�=�ϙ�ju�������G�玗g��s���Ɠ��m�W����V,ltӯ�=R�0|=.Q�#
�Ҝ������w.��:�dL����@g�q��2�F�9˝��� �R�����|@��g�
��o ͒�=�
5�}���ͪݱ�� �I��p��^�Um�*@��|��^&y{*���x��s�BZ���`�n�וm*;d!�16�&��� n{��� �LX��w���ܼH�is���z����4�5��WI�̢�3����i[x��7����ɵa����q���։0�}�� f�]J�������X"u}�g������A�lĖ��_Z@��� Ҕ)8R�Q��|���c	�ݕ0��C��: �I[�U�RË��G����%W����B�ҊV;�U n,!���8��@��K| �]�f^���5��ii�(�D��A�����a)���K�$�O	u�R(���8�<�ɹd�u�M���O22����"�dz�����1���"�ߗ^�S�]�o���ұ��(��G�k, �6S2Xݯ{wn9d&%p��n�O5P��;>�-��^�|�d�y�L�FZ3l�jd�0�k`\r�/�@?p@�����h�I�y3+��sY��$�^҈�����DعV�ǵ
3�R�!KMt.���X���Ыӫ<5�d�sjyy ��	s�P�h@��P�۩Pfb%Z4��Ы�����7�o��;�,C���S�j��܂,�U�k>ߑ8}�)�c�\�E�e過���l˨/�ۜ���C�&C�H�΀nA����;��=��Ғ'���b��{�Fki��z�ú�u��Sg̻�瘷f��g�r�݅+{V��t�a��H+�ޠض�oq��?� N��Y-o͏?�߻2�MC���~�jA�c �՛�@<h#�q�T��2D����Y)˷��;�a_@0Vnl��(�\���&EśxT�*b7�Å����|�-�`�0�~9�|���x�������m,l��-,���;ɩ2�A@�C�F��hM��t8�0Rd?��Ί�L��hSw��Q�i� �|�\��0�}Z��z$�6�{B�@�`�)�����y
�F[\I����'/^�>�Q��ح�a�vXI��N��-�*}�
+���y0� œh�)h�(���Zw�(���ʾ͎��1��]�`Y\?�9F
�Ki>@��_�Qu���]�n@�C��xX*���b�sB�1������E9*9 b���7�Pb�Ҡý��2߱�+b]�ݚ��V�hLc��$.��ho�*�)�Z�e����K�l߿�#��OaC��p��I��J��`/R���i��z����n�R�Cd�2�:�>F��j�_��jk���]����?QzQ/)f�����LL�q�-�/��n�������A^&���p:���׼o��(���\Z�.}��i�R_O�U�>��/5�y�Dd�2*��/C��sn�DS���`E
���I02���_�TT����0a���V:�ƚ��z�e��(�5 %���Z�k4ߊ8��%$E��9Q�،��h�8 :۬Q�w#+�5�X�������ڴU���߉�㱪EY�����n�cz
�"�;�r_U�ş�lC���+��l��Y<?ޫB��m��|���M�4�����GHu����F����U(Cu�����<��V�kP�7�ͷN�q�s��Lt�	5n���s���U�X7e|�����뾯?n[9�0炷+��e���,��l^#�}5�JV7�J���y���^���W��(��#486�;�"��"����M����Ƴ���%�Z`��D�K���(q�:GK�]��\��3�U����6c�o�-��4 ���PK���`��!GxU��tzf;u��R���Z�������*�!�N%?�R��+�UT�XYx��p�7�U&��-�Q=���Ԍ�Fy��y�OA�B	(U��@nt�u�FrK�u��
gl)r�Xl�ר�m3;h�����Z$i��ߒ�>[�Ci��:�9L�ޞT�(U$Hӊ2*��R��n�Co{K����s��%3t�X�dź7����(H�[bDI���Y)�o�G�,���g:"����Ɏ�2[tm;ʽ��/��!� �=�v���؏��	cov���_-x{��!�^�+�oV:9;�0���-���u�1�=1~��7$B�.�02$�����ŕt���3b��R^6eriU�E/�_L�1�Ǵ]Dip�&(�3�o�I@V7�
��K�fH%�&�|���i?^VX]��I��;Tr��S~D���a I�"
 ��.����4Nw��@Bӻ�W�s��lE�P=mL� ;;#�?}+��Iq_[ ����N�ze͖d��7�Ǽ#we��Q��5F8��6Č��������(�]}}��p+ʠX�xX2���E�����R�O��e�T1�=�y�] џ\\lQHy,�sM�WX�T='��EUN�8`'���6�ԣۖ281��^"	��]ҶB�:��S��������'�h�E���'�j|�̣�%���y��ci�(��W�a'��$A��^���M꿵>[�)*0;�y��Z�p^�7��g���5�9_�ǔ�w��\E� ώ��\���dZ�G���+z��9S��Y�lC+*^�Γ T��j���~0�}�s7���:B!��4X ����{ٗ�v���h�c��ݝ�����%ø�o�iD���5/­�Ԝ9��0�ϋޞ����hЕ)��3���q��@:��\ސ�3I��Yo��˃!01�
�M�Y�k�:׮���f� {�;��r;��qjq�ы|1�S1m�
C�B����{�<�}b���|R����qV	3�`����$L��.# �@4���`K��\��M�P3����F�6'qm��M,�����zy���8�k?�د;^�e[h��*i�1f�5��ٓ�%뚅0�м�?4���}��}nW��k�4^J���ey�����bA�c��&�&�H��bThD��~3�V���o&�G�PZs��t[*=�u����"���R�4�iSӴ��ز���XK�!߶�=�v:y�@�(e�(d�z1 ĴΫ��(������|�WVL&�7��.ۤĩHW7��gMe-�c�*��m�?	f`er-Pq��6����b�ZH˅(Ӈz��*����j���Nъ�y
��<\Q�U�I����u��xH7q����/��0����6x�d��`�47��'�����T��E�ة�V)͑�̣�����-p>9�ʏw��K�Ph:�h1���9j�4$K��[VV����r����Y0�����c�&���-������6b�'��Ƌ��L
�+h@$��o�6N����Xb��Y��������5�E�BEjm$�����}8i����P6S5ï����8���jv�c0_�D�6Xk�*��T�r9���e8Y��cAΡ�ژ+w�ɉYW�9��Y��5Z�U�ӣ�7=�	��!A����ðj&�X��W���s�#b�S(�Y�j}~��"�䐓^�7��I��PmY8�C��߭�:z��=]=D�w]�����/�-���I�E�CmF]���_��/���A�4Ma�Q~L�r�aR����D(^��|�[:q!݆��T�8K�{Lq�6v�[h��Xtt�5,�+�]��1��G������]�r��c� %Ȭ�Lv������o�po�ꗨ'4�����j��ן���Ԋ�Mg�H�6z����NybY'��`(����)u��ٜ�'`8�Ÿ�1Ԕ���.�J�~*���Sh(�ދ\H}X��*�G&��10�-wl��hvp�Y�>��c����UaGd�$�qJ�'?���@Ӯ]r9�5!�o��ϦT7�=�����z�	r´���~,�'4�q�6DG5��*郙�$Ba!(_�QY�"����*y��Sb]��BлR]n�~�O�+���W7�?g�iMK��x��{ވeNJ��yQ���McMÔV����#D�^
�W����]��瘎:����������קW^�
\�h�>�.��^��>��I���%�)�ݟ4�e?��h�TB���%������<v�LI���?m�%)Sa��qUP��>�\}.�uhZ����9LܜLf]Ȣ�%�#aꭧ=�9їZ7"�Ay&5�l��h���O\�տ�yy�c(��x�E>�"R��d�m�Q�
fE�r̸�]0��Xq�18�71ū�d�EЏ� ?�������#��0���,�Q�d��BJ��:��`X��Ջby* ��d@!��m=]�*�ZD��6
ϯ�����K��"lL͚��H+�ӹc�oz��-����� �GN�|�8��#0i��_1���U��yb@ +R�+3��A���ҝ�I�����x��*���%��(�:�9�L��ӗt��#�0ݧмZ��x�!if��رŜ�y�l�����,�<вR���\R8�Q��>����yłS��c��4�o������m~4�h���	��=&s�/h��pI>���b:;�h02*?M-����0�6	h��Zb�u��S�u^��Y�f]�Gbd &��R����Y�4�)0
���2���C��O�r��o4, b�o��v%�B�f,K��I"OWWE	R�9_�x茂����E�η&�g�� ;1�R���ˑ@%>�jp�H �X��}j�d��<�س�2O��	»6E��z�2��������\>q���.t�����C[p�Mr��rk�\0�
A��}�=K�ݮ��q}��ɟ�fe���-��&�
~���*`e�5O�Su�$x�/��=�͕��υ��hA��� �{T�{�-�8���h%���C�B6;K<ڇ7#%ƕ�!U�\��ONP�.��#&���Vb�5҈�
C���G���*�m���'���X�/�J[�Y�De��=����+���u:K2T}�����*�պ}���Z�����Kϑ��X���1�=����_z��>�\�*K:D�5�ڡ�����C�U�0� c�e�g�b��0J�AΏA��gz����V��^�0�o�J2+���Y�:����	����B��G�1��Q�?��r�\,��uƢo6Y�c<*@���N�ޓ6R��\�k��_�����=��d������t'eA���U�z�nGn�h����&���S�~>	���+U�i��·R����
����������>�,�n��-*�>:,m�/��6m����n��Ǫ�hu�g���E��SQX1��F��<�$	#%D�Pv\T+vGh�����x�T�W.u��Tts�I�u��V�Ut������g'_ޟ�����?�`��݁1�j0*����t�o�H���8_�d$���81� mQ`�;/}�Nr��L�x����G�������� �<��$ 
KK�g�^�W�}�xq�RЅS���|��[���Jށˢ�\(��?�&�;<-,��d�{�wC���V-x�C�Kzb`(���\`)/�6]���0�8)�1- s��
�x��'�XJ4�M�SkZ%bR���Z8̒&��?T����Dɂ���}/ܽ��-D7,��d_�H�Ǜ���P�D������:�): �Ϸ��t�z����1-�MH�*ư`KN'�����&�ɡ^3�7�3y�!J��j,����kbh���H'y0JJմ���4�X�?����#S��Eu2�l�J� ��N�$P�,�ۋO��nL��}�|���4�ݮ-�ދ��f�g��.L�a�e⯂��6]IP����g���k
�d2�U2Fl��Ζ��>JNta�'�a��zH�bQ�cT_\�T�j�y�!	�FG�_[ج#>$FY10��Lن/g���]���5q�,�u
��~�t�������o�z��e����ԉ^\^��ެ�{Q����5Ŋ��o�YP�u�D�25��4��40��x>��\��cĪ�q���/��2�����[��;,�$j7���a�t �g�E�~Ʌ�C�Z�*k�����g���A$j�C��b�Rc
����g%���	=4oz6+����t�N={��;�im�6��|�m��ɤ9菊���m�!�O1P˪�� b��滫is����@c��2)��B|8�+�%�ͥJ�Z-�����������If��Tı=����'ܩiX!CT��2�H�p;H3sP����秘	��ry�����@�+ȡ������|t����b�+�_�k@U��������T`��G�������1M��A2*{�]�v�&dq�=ޏ��]��t��� �|�W(�'�z/j��[?>�����%@U��AI�2 ��"Ud&cN��x	X�������8�r�v^�Q4�ʞ���ק t`����"���W����u���s�l.p3|�����o�\�˷��x������������(W��5I�Q�k�GLG%���C嬱d�pB�����d��l����W��{x�g{b����F)&��%F����ui�V`��"����	};��H��{J _E�>���l|��b��1�x!���X�w���P�����9�ǈ��OA������y/ ^��*ζ�&�Ǿ;����
̈xd{
��?Z���O���O.�{T-E����#��Y��{�m�ݍsz���~��bCn9x?�P��sOu͚ӑ�q^'���z�� �b-��;mz�1����I�	�'ḥ����sKv����OqB����Ƿ�5�Vi�'�Fp֚����GH�$���ӹ^��������9)��f���zK��Wi�aN��xѥM�����k���>��>�2eL�hڐ��չ��nVAT�'�2��m47s
�잡!�p]��F�{K���XH��0msdjp]x���.�Y7���G[�C�b��aP�9�5 �-�\��Nw�Y��#�b�;H�W�'��>�Z�P�"�̓�#��E)pez�k�"A� 3���v�G��Ds[��l|P�4�#͚G��0T�g:H7g�h�)hY��nك��� qć��8�ι��Wj~�ʽ0�\�`X6q_Lz� ս5��R���5��l���_��Ά��Z�v��EJ�����[��"�0Ҋ*^��:�K�{\�Ǆ���$��~��i�r*�9Z����X��o��c��ѧ�L��¡�g!Гw�H]�������
(����-Ӟ���~",]��`��mW�3T���;.�����u_`^x:��3���P1g�ϸd��l�A9Ǻ�~�՜<6z�����^쾉�(㉲fd�����Q�iZ�x�`����M	��EF�	����og�Tiw_�B��W�)�jhP
�+�ml�t���)>����U��2��;��n*���[dkÏ�&��~�*�DIcW��_#���壏�M8P8ԾBzϱ�ƈm]b>Ƀ)���2D�<�$'?1=8ɂ�����Ϙ�ޣ���=���qZ���> g]��Y�?հ?K����W;��2$��C���bQ�IkX��mxƍ�c?]7G8�$dS�- ��lK�IpH����i�x��J7�y��m��d9�����vȢ;.`�]^���T񂝜�yt�������<J�'�8?~��V�i\��t���x<�˅�i��������r�l�	$P~YE�^����`�&7�0�V�"�y��0'ƫ"�����o��h7�՚��
��k�H�By8=�����O'�O�\�ʌ�v�oo1�*)H�h�� ���ǰ_��>�Ҥ�'���4d�:6�{�͡�7�!A�A<�K[?ȣ* ��T��B�����
��֬g��ez���)��75�[ĩ>ム�r%v<s'���U�x�ҷWB��?��˝:d�b��/�콪x&{�\�RC�b5m���i���@39*�[���"T�o3!�zo��;Sq�q�8y"�l7��\)0�&�ꊽGh�V��7� ׳kЊ�.�ٔE��ҫ�F�7H��>�,��V�FZ��k��HӔ�;��ǡ>Q�7>w��l��{���|��
�G�//�(#	 ��
�P�U�L�;a�'���рb����:!��]t]r�D��Q5i��wE���d4�:7h�^�ш�/wk"2��i�/����E��{�[�\DЎ����ύ9���N�=��ߕ�	��02_*��(�6WGh$���*��(��Ӟ�}�,g j�� �Z��\�O��]/�K�38���GF�G(n}@BH�wQmk�W��%��Ikx �s�X7>���
a��l���->!��B(�k�3� ����k���]���YC�p���G��c^2p��!�贆�]��G�.JZ'��U�B�V� I��(LP����Ȉ�wU+q[c���>�a��>�9[��v�ր�!�BG�x��o���k���}�i�
�Mx�����c�i�z�O7���+ײ�IS��*?l�u	�W4�`�"$�KN�}���zW�i~�@���)�r��
�J�M�-S���s(ǸF��{.�k�� �3Br`/�4��p���>��M1��J	��>�F�F~�~�C�ù��D�,�?�.���X�e;'>�x�3w��t�6��'�Z��ĻI�(m8�dM�hxAǻ(�}�Yyq�X;k~0��3D��'Z��k��6�\2.5ސ�Q��Y�� ,�;����,�C����Y�Y�-�5Kb����NG�7S
�~�[d�j�BM���P�2���*<|�?[vӾ�����c���}�sq�qق��dx4�+ჾ������ܴX��ڦ�J2���#��\�/��!����v�
���CY�;T�C��
�Y�
�;u�IDp�֞C��cԜ�Y��z��A���ư�a��"�N�t�#3�oV�D�_��ݏ����ra{��),�8o�r��8���SзR��q�� *(Ъ;�M�7�?��"��R��i�lsgӑ��E���S�Da�i��ԋ����W���V�Zw�@��(�X$�=>�*��H��޸����^��6p�����od�{�_
��O*l'i�υ�Q���B�3	Yi�C��Y�kͶR����v+`��A�r��+5Lo���%?o|E�92��B�����)�R!�/LGC<��=����<WVg�`q�I�����a�SÂ��KX��6¯���5^�R��{O�Z�T��SRjR@֍�F��R���G?����p'��bf���|�����>� �z�s�AomqM2`�\����S8�SȨg��`������2{�Q��
>D�ȴ�4bQ x�h���FÆ�
��j	PixQ�;&E��V_�� �%GN��ꥬ�z�ӯ�
�]�Tv;�d�D��S.-[)� 	������}+�3������{s+�~�~|�ܲ�}��L�������8��tTՕ4E� ��3���F���?�/����G�-g�p�:����.xFC��� X�'4�P�r���I��2�����p�QƑj�ftmp����䟖�A<�ITg�ɔ��ŽBnԇ��t��� k���I���Q��R���Ř�u����ӎw�� tXfj-Y�5��|�ॢ�F�/��A�Lis� ��;��"�����<R|���9���t���0���eHע�eG�!A�Bk��������Qdp�[=L�;�+r%<�܂ H�QP���(&>� ׼���i��U��N2T2o]}��4�w�~���S�{��7�a�hU�0���yx�� \N.�}/�;�媧;�8B��(`���$`��@�v٦�4���h ��w"�VTż��� �S��p�POF�����rέ��4X���*zp��<�B���AUo�҆�/��ݪ�W>:m�tN�"��?�i�]�� ����|f��q��(O\��b�����[�ԋ٧sR>V�n��b�|3�/}���4
w����'����vsk6v˓�DְE���@�f����Dà��
|a��M��̺��q�,;�r5�>�ؽ!R<�$��u�w nהb�Wm�O�w<���������f*�O��bZ�� ���7���ML����+��js���J��K�x@�f��T O�)`�7x�8.!��8n�7�� ��K��L�p������0��,b��a޵��~�������}�!A��>v2k�a��S�y�-�\ ��"}�y�ߣ+��0>�f��*0#0�8�:�
�EW�u-Ƀv��-f��R�Gf@@��,��5l�r�6���F�2�Fz������K��|j!"�P)ʲ�r YF��yW�Z��ᴯ���I"�܅Н[oX\Xǎ�~����{i;K.�;e�QͲrɈ��~��
Anzғ�����v�x6��ST�&vW�fd�j���Yq�KyE�y�K���)����Ycr�H��������� �2%��s�sk�Q�K��	�>�'�HV� ��K ��U�����N荽?�_ �J
m�ԕ�: T�5!��dK��F/��v����#�<&Ӟ�"z������\:�g��4�Rt�01.|̠��҉!� ���А���v��w�⇔�5:M׸m̷vP�A	�2! �s3*��8iq[sz�y�DU=@�P�6?8@�6�/kb��lwY��?�x����Jb�˶#�]j3:{�(�BJF7ۄrxb�ߖi�U6�^hc�b�6�$�h�8�/��Y3�����l��Z>�?��OW[N`���P��J�B��0�� B@�.P9s:FB.�ns94�?N �k,�Ӂp��y��	��l�+8	g�d���`�J~�'x���9���pT�JGB���K_&^��x�Cj�3P?�U[�� ֪�������2L���7�$x��FB��_H�}.��mB�f݃�p�Q"�܉5���5XE��'4�7����/���ć@ y͜��E&��d��Ib�Q����B�;��f���B
��g���wmD��蹰��R�HR�<�ƛ��c��I�aZbh�P����G/����^�>���Y�� #ʧD�s7�P���G6S(����KUB���L�3���L� �*)/94J����@*o�z����;)�	2���cݐ�d\�g����/�h�����������|����ܶ�ھq鯘!��E�&�}�a���-'�f7� U7��2G���Y�9����o%Ȳ_VA�&T��׌ ���b�ӽV��H㧶d>jl2�i����+��$�Z��W:�����9k�B����Ҩ�LH������ÖL�].:��ИƔ��oG�"���B
`,��}t7����D`l?�f}����D�X�Tk���Ĩ
dC�>k�%��4�u�|�(C����tz�O�[���	�p/[ r{�Օ{�|�������X��(��Q�4C6 u>��nvr�1�y����![���&n+0��Œ�d��Y_&�ڍ�X[%�!Rwߍ>C��=4����
�
iO9�;�v������Kmė���p���$�(Ftdb3��p��>����$����)F~�Y��d"�{_�躳.ss��uqS�2�3pW�0,�d>!��\X��U��qB�K��&Ĕ
����]eq�wg�P\�c�Co_�6N��<�-�
�r]i����ɩG��	=��=��%��.���!@�;i*��r��� $f\"��9���&Y���� Qg0x9B*�)t#��w��������%���i?Ѕ�eTMN|�u�jj2J;��|ms����n?�=� R�B�:��v��/&q!�D�=3(VP�=RM��Gbq�߄�V�[�7k�L}I�ߩ�"�����5�MN3=�)ɜ��t��p^��ek}&�k=ެ;U���*�;��&�M��5�>ެf�����z�X�!�p����~ϳ|�¶#}�C�0Z��B)��x�k���#
Bi�^�A���c%;��aK+\�����Ʒ������/�A��������JD���/P�ȢqC����L\���\F§��\�),j�]��Pu�>�T^�+2���U���`�=%�W���K ���ڪq�����A!��M/�	�_Fe��l
��ӸF��`�R�N�J�e�y��<B��̞�=�e?��@~&$�U*VBl� ��X��Z�T"R���p��ewO]p}�_
��L�H4�-7�T��N�n�t�/�Pr(�ĐϔR�hY��U�Uv���N�i�B�+a�~Q��k1���ކh#�_������fEPy�Ua����T�d�QY������{�����p;�s����>��ņ_`#�2�ܜ�N����Gџ�b}���\�k��H��1okuP�|�I[f@��ӷ��p�i�="�!������U|^Z4Ά7��;ԁ�?�ғ�ā�s6��y@d_��O��t�*}zZT��-�����:(�o�CC���Z_NccN����+Ǯ/>UȲ;��ӂD@%Zdc�h�H3gW��4��%q�._l���#9��=���<�N0��K�W7��QF/�(1�C�@M�h�uh����\��J���1L�幊P��(g����O������d�ӴoI��O?FPW�����x"��]pc?����u���r�莼��B吉#٨8�{P>���ֽ��z�.��׏B���Y�����MYռn��T8)����	˼$yL���WY��i.�#��[��V �D��:�\u��@h��߷��Ξ]��K�T���s�hT �����֩��.���g���Ŭ�h����p^.��B����\~ۙ�Ih�D���2�^���D� �� ��=�TKB�Q����-ŶEFK�1]�x���&��Q��S��j��и�Ԝ蹜�9���5���+����J�2$��t �͏gM,�?�����{⛚u��:ۇ��I[l�h��?��p�������ҡ��-���3� N4c;��E#L��%}fV���| c1J�7�2A�*����L.c�_y��L2�� YP>tġ���dr>M���ӹ4B!z��|6(��lB�O�>�W�Ys��2�{�Q��@�4oE���a��dH��}���e��	bh�)Ƥ�	��&b�nQ������#�����X�H��cl���2 +(���M�̌��I�0qv���ވ���&�G��K�b����*:���D�<�Ѣ���߈$����z�қ0�H�Xs	��?��92&�E�o|�@�) )&=4�R&"a_�8�0�����pBpN�K�SY�U�a��Q�X�T�W0wI���u�05WT����_��WG�¾��7�3*�v��?��˄��R��}���R���w,c2��ض��"��D)%�Ъ_���h�Qkkb����r���.��aĂ(����R��6/Y��by;�lp�ԛ��"��~�A����ջ2��ٱ�&ja��u���:�I�VwMh�{�[�	!L�yv\	�P{J'��`��_tO��@���k�6���V�RK��+�Ǎ)�:���l��~������;*	��P�� 2'��S����*X3�`�1(��2���3��X�~��[�W<��1�$"xQ+$�AJ�̫��y`�K�6a/�VKf����h�V�&$��LȌ��,�G�=�˯�pDÎ�e_�����*�^�k9�|�N�'�����_�R�r]@�ͦ�P\���^�/�d-�B��x�T�m���[�i���x����y�^h��M��@ؾ��X��g@R���SWc�B�����8�F&�}@7��7j�7��ZĈ��
�w,S�W��=�����q�ya"`�v��6�������9���d���3�0M�Ǳ�l~��e�ޮ�Ue��������Y��A�P{���8M(5�e��zS�i���Ԭ]���b`�ݜSf�H?�60��v{�݀�r�ѹj4}�EwqeS�s�ro}��/����:p��L�$ʙ�����.ߙ� �/T��ɥ(��8�g�4���$�w�p�K�4�^�����|��S����KqL��>���|�S`����g���X�̚�o<���ͫ�`m~�d�;������uFu��a�k<9OuZ�%���ꉗ���%)9Ȓ����A��]Q�Rs��vJ��E�q�V���q��ڋ��LH����W7�{�M��4��K�bt�	Ϳi�X/.����1`�P�!���cL6O>���bc����ԗ��Ud*7����><x$hƫ}@?ǍU�������g@�(ңοb6���{@%��I�Ǐ�pk�(�%��btJ����i�[��)ݢ����r��]�B���WY��_P 
�UdKp��rC�I=+J�t�>)/R�^�/�q�>Y�m��X& �!��~T����.?	�ҟ'�QklzA�ΞF[�Pj#���ҥ��[U��v��[95��J��*�̨����o�}�|�,~�<�����8 ����`���A��Ýl\cٕ�s=��7�	�)E�09}>�����0h�vv�dX���S�}tp�bi�B�2�ŀ���!�ȍ��\��E�m3jǊ��4�͕}�DF<�Z� ���x����n�����J�r��F�"1t�hcd�3�Ձ����2���{���)9L����pU�{��3����Kb��w���>5����n�J�(k�����c���X-�2[S�R6����~���Ǆr]����G�X4���C27��$Y׭M .W�Ir���j�'��"��hG�leXe����nHt��$��L����'�C�(��G��١�R6���}V����(��%@�\�2�X��I��gB�Ln'�U`Xi�Suo��@��ߤvb���#BhU�8�����0a�ƙ���=�[\�T��U��p��,#��f�G9��ң@�	Ď��H��k�~�E���oKqL�M�f¥�� W�l �����=Y��s�Y*��
��R��:gع��� �*K�{�j��5߷�7g�tXwvcz˛���x����OX�3��^FFD�Sî#�G���4��p�}�X���f=����T�A�~�J(������_v櫴�ͤ wu�P�''ay����-^�����$�����ߚ�v����;��4�sm����}{W���*����	�;�΄�i<joai�:;A��Q�q�� -m����h�N��4�^��*�@���08�Pa��,���QxFMQ����!�Ͳ��\�w��$������f����J;.�o1X�c�G����8�~��P8шWgJ�=_S��h<���	(�?�p�������;��N�?�_�������=�� t{�q�OjO�XQ��t~�/�^���j�2�_V~Eʲ�A;Q�,V��7�zA�Q��������#WI�&~mz&�S�2=��~�uyi~T�@,F��ܞ�bJn[�I�95 ��"]Q��J��YY���g��?V�j�#�.��Bn�$c�y���p����w���̚m��O�
]�_Rt�5��o4)���&��˂c���>�yu�	
h�����4�8�D�(o�lx�y����X��L�ht�r[8Li�t��6��'D��Qr)��
����1o=U��!�
X �G����OL�0�)@��,��Je�I�t�v�r苪.D#�����N�m!��9��"6h%X5�=	Е��!�{�=~�>ˤMH'%J������K*�L�7;����d!kt�� I
�.�உR}]�z<��)As���x���m��n0&!Y�n%��1�XI�}"_���K�Ǐ��<���;z͓�T� l��H[��NC�Y�i���B�W!����ƀ5��7�J�~�R �z=��(��O��V'��fVכ"m�/u�n��(P&�ϖ�;�V�����N$�M�����\�b�����{hh��"3��0�!�<T�I}s��q{�yaUr0��b &WX葋�쩐�T�|�J�Ö1���)�?P�6��oQ������Oy�`�2������5�B�EY����u��'c�Pm������ɦV���k�v�yN�iv�\0o'�dV ��A�ѿ���y�S���C�F^�'"���}�?�jEa��ڑ����h��T̑2�տ����|	]��R����W�ı�-'�����x_��!�[�=ՂAa7?�*+J`��1Sk�f�8��@�I�ԥ�l�q��J�/��$��]*{�#���ٓ��dy��i�D�i�WH�n5��;�A�C�����U�ٜ�A�o�H��R�3�,�v01�/�2fj�,�J��"6mH�LZ'����SiO,�	+`�W\;24j?��j�}?/���q��P�s{6I3����ph��$A�����ƶ�����"!(,@����Q������^�'{vE1(9 �׌6�}l�r"���X�MO��	Ѻ�ñu�Nsb
['�{c������lH��y��s
;p��bO�k�\V|���,x������,�� �>o����g�c�5��0&\��y��V8�~�Q2����$^Җ�j��"B�~q��QԪ�.0��_EO���� �fD�LE�&&g ��~�,��,\�H�4���w�h˕cf�.�(�P��?�h�Dع�hu�zi�Aϒ�_lfxؤq4a�����%.�`����2Ç.�Nw7ɗ[I����E�-���}oOF���b�BHW7Z�c;���f��}M�"i��o�{���S�,Q���|M:��0̓���<��-��=� V,��-�c���-gV����Zcܺ@:��kJU1��� +
��"���In�
[9�e��Vp:3�Q�{b���r�'񿵩ʥX��\5��6Q	����R�.JƠl-���E4qV�t�8��1���g"U�.�UwG��{�
t"��Yx�S�#�T�	Q�������s��	���N�L�ĥ�7�n۷����,m�p��Cs�21,f�C�讁�*g��)8�1�OVb��x���:x�<>��|O]%[�:gt.#����N�_�` e�+Ш����ݿ���S��s7C5MQ?�K{��jd.�p�j/�%�g�a�]���W��]7is�۾����:�n��\���j���"��yP�?�..&�	=��qPi{�
���4���j�����>�_K@q����~tטB����Q�0!z�9���ތ'.�yғ���7U�{I1���+ٝ��u�c��5� ����WP��1���]�����WI:��x��<ԓ�hnOȭ��KW���\ p�i���d@9��u��Fq������BCn�Z8h���OT�?�Mz֕��>bU����+�W|�";iƫLJ����n�-`�7�MBE��O�S�� ���R�#2�i@ I�gVP�#M!��xi�^ߨ-����u
�t}� u3iޡ>ps�]�3�kj�-�뎝���7���Q ��]��2�0h�V�]�x�&��;GndO͵ًq�����*��Mw���M�Ƴ�~��kr�$�:ɕ��a���%�4��r�6�y6%*/�n�>�ᤇ�f9
Ԯ� �M3�q*�a��p?(�����g��Id9mE��۰���!F�*[џ�qH�Q�o�Y��X֊�H�VM,�9��s4���	K�'�Լr�C��{���E���^�(c�s������^֖����
,�-1���z���W��Ӝ�m_��2�NU�<��y����"�HhM澏�xT)%��45?�:��s���ZQ,��8���&�Sۖi��E�09Kcg}��\�����I�;�ǩ��U�`���gH�ڂ��~4L?��(�ؼC��� q�T��`��(��C�L�-����+�!�F�w�"��u�}�g�5Ŕ!$���#�J���o~8��3�r�ǟm�FV^ut��'澿i/���`^��Ҵd���Vd�����l5���<%
��h)p��5��}f�r����:FR��ɜt�\�m/+����.�'�xi16&y-Z��HLi-��<�e��@������{���ߙ�Ė��K��)r�d�V�wY',�(K���=]�&gxr<����y��i{9�x�M&�^c�����I�j����y� c�3W�_�חK@׹�8��D�̥�N];�Ł삡�9G��B�$V���e�y�&�v:�<<�ՠ����0�m�upA�=��(|���
�v��]�0��G~N��Gg��U�˨�0���.�u��]e_��܋9|�>=<�ߊ:�_�O+J��@���85�`BCZ�;�ൌ��5�{�����&1JZ'�8��$���_ω��)ڠ�_d�M�|�(�<�����J���\�x�/$Bۇ\�m���Q��˝�r0q�&C^�k�vc@T~�������,�1'r+GE뢏m0��qx��Y[�u\�7æ^�8�M2��PS���}�����ݸ���f�-����cQ��J�Gy�Ks��ğ����߼M��q�2)�t�u<	?P�^�<&�Kh�����T]1@=�>y�� ��Mm"-뢹�d�������HR���r����#��F��M����F���_"}x���)��e���Z8.Ha5G�b�����r���bo"5�FȄp�(�I�߰ЃBUp�"F=�����}V
��t�|� Qb.�����Z�1;���߭�3-i|=Z�۫la�1Pq�����=\ �J�n1���
hD��M�c
=��nI.*����%��cePIC0�8 ����r�~*H��'l�v�N��������/�&rs��p::��=\��`�Hb�Mo��*�5�[p#��4?C�G���pVBALV���	Xu�*  �i�hg^ؕ'�üN�	G�0�6E&%o\E]l�������.����<��g`�%������H2-3��Q+��;�^��x�L�����J�%��)�V�,�C}�9�I��yW���é��Ku�
e��m��R�^��p��} G�N����1 ���[Y���)^+s�RF�w��;m��{1���	e��Q�n3O�#}��
\�/���u�h-��VU�~ϑv����Dp\�; ̊H�S������Lz��Cʽ-��`��\�J��j���앋�qT͗�����$�䔁FC=��%�6_�jع�7�d��*��HG��ճw8���!�zjQ.|�"�~�����Y�vG#�n.�q+���կ���m�/G��D���F aV�r�4r��<��~K_�H�&�WX��n���mG�A���f�DE���*�����o�ff��V�:T�ئ�?]qNr��a���ӻ�ʹqtbg�����fP��xpIɇ�м����U�9C�(0߬SGS6z���7�r2�F�܌\�s�����P|��&�d�t��!t��ql����2����*/�Ǫ{���׈�3t�ko�a�����k._�������|)��&ʫ��umK��̶'9�7�k�1����r��'���δ�
�Biw�� ���Dh�8�$N��u�Nx�b�c`�7�V��	�W��:ĺc��-�(͖D\�QѻB�6�[�4�'{�����4�6ʙ��g?`�����}*I���=��T�����g������;X����(��Ns�.�@��ٳC��6A��u�|y�@:gH���m�����1���AH֌�x�������SP-���@����<����,
�/�z;�~E��ő�$�N>�d�������b�1-�����Y
:r�+���}�ذi1��� C���c9��V����׭jJ�!�C^���`����[�����<��\���`��x;*=	�\��`��.�__�P��	1���y*��7q,4M �@8�v_0;ii��Ul�$c����,*��;IYs,N߸j�����ް`op���س%jIԆS�t�'��im�L�>�s_��=�-o���o�H�7\���,#��Gq���a��XCT�*|9Ri��~k`����*/�o	��R�[���b:GX�>!�8���a�Cf@xKs��� �_���.^nSP���"�2��\�R�%�W���f�w�ժ��N1�U�w�Sq"�D�۴\EĖ*D���칺��x����L�{�M�[}Eоࡵo.�ӼZ�*ڀ�A�H�ΟO��X��K �����0�c�Y5�L����(�G��2e�(bv����9C�Ҷ3�³ޔ���M�'�Y ��ۆ W<�#��B�H7vf��6ٱ��EM�V�R�mG�c���?><�N�g���Q�n��<�������!�7���5E���hp��o%�^��L{�\������:XM��.�8�i�7k��ϴ����]���b�YTg�`�[�T��6a�E��Âq��)���c@��-��/ēC�l���������	Q@��vw�R��-�Ta����o�c�����._wƶ>`��m���k������r:�:�K� 	�TKU»�.������V�Ks@ Uuf#�-��!���B,�����CX��!%w�*s��Jd.U-��%��R�t5��^��;��������t|�/�L��H�ވ�L&vUb�������f��0�/�,�Oۓ��+�����ԫH�����G3˧�`�&76�]&sہ��%`gI{���#,ڸ�h���2�������@uj[���%�_(d���&�r��Pz^��
S��h[��O	�̇L�f=OL��Mۼ�"ƷIc����"6�p�{ߜ�$���	Q��4G�F����pd>���JģZr6VYL5��3d�t�O9�
+�x�� -�:=�����5�W�!`^����^����R�z?�
�N�>��p���� %~?/��>X�WĬ{����ѡ�Jm+�85�g�n�\�,q�UG]޻�
��p��c=-^"b�������7v��ziM���O��/�@9߿	U�����g8�7>����S�	����ݜ�~h1|��-(ƾ~]��
r��-c�"Pm�򘚮��6�B8���- ��L�3��4@��B"�kf�sR�����?>�a[q�¯;g�7�;�� ��-�z]3��0�Dg���l5}9>ǃO �⽂{�H�YԱ�˹�*�b�Ք@��a��g$����g]���ĝ�@n�M�����e�?i�v��]�3��t��:N� �68P��)�_x-a�hޜ��'����E2F����)êּ�}J�L6i(���Y��gkF{F��|]<��j��6P¢���Tc�[����C�Ҧ	9Yܼ�t�f�[�PWq�� �?��U�́�܈��e��_���f"3������]]�JD=gMHE���(�D��SY�bZ^P�ˬĖ�����W��w���V�J�?��cy��Es�\$t�:��$����oOLR���6���������VjBRv�wg�8Q������(X�����T+���l����i	1��z�P���W1�Û�-2�3�J|�_�gǮ��Vuw��f54�ctb��q�T��e�̖|R*�����9n�D(+�_@�>vø��f�X�����4E�s3
���<3Ո�g���5�W�(�iJA��_w �:1�.ܬ�k<e���S��J8���(�7zP	����+W:d�.us*^O#�}l�ga��4�a^_����˖ J�^��`�W�I`�ϡW�:&FN@'1��si�������"�ҫK��+�^y�^�pk͍�?��͠���{��&��y�7cS��LI�O��W~/7����\F���R� 0?�[; ���T�+¦�0y�[���`�����������䲴�]A�OZm�dF��8��>���p=}dZ2������l�DG�,$��}/�e%=���v�Ѯ[IW���Pjv������$����i�Dr��~�l����T��{ŁI̹�/��!�J�>W�] `����q�5È6KNu�
��N�������i�z�3:�5*-�<���36��fӿ�5�T��8��P���0|��1���.�=*�2�v�9�{�����{7��V��~�.�8f��Rjf���iz_��@�"�aF?����p�����?Ü��3HJ�Y�O�+���㕕\X����6�CƑ�#�&��ʊ�h'P��rET;�E�����ZO3��r��^����cT���+_8��'LJ���3F<��[�� W\���:�1ݡ�CM�Z]&�kvy�VV�ڂ�,��7��@,�W��N�pq�`}rȍ>�E��W@������E�H�,�`�M{S�+5	��?B��l2����Hw����,I5!�wu,!BKV�\��`�nx]�#�T�!�}[Ӱ���c�O$`2M���=�,�&�㵦Γ���6�Z��0h3��TR�x��d�+�?S(d�g��9p�-<5��$��C��W{��N�4jYfpY�]Be\?&���)Yn+����帉��IkU�JRC�t��^� .��W�_��Yd�k��{�?��5�ri`QO�$Urz�rD�(-���p1�'m�CB��n6���;��+��
k��{_ч~�t9A�m��QO&�j�,P�kςV����S��*��	}=u�C?�V'gj�7{�G��j�����v(������ا�=?�<'��d�E��=�}Y�sn�$;����7�־�E�'�M^�#���/V3㞎=&ȍ=�%/I >z�X��z�m�A�4,?E��������f��x{e<�1G��ĉ���wtQ���^10�������mdo<S�ԐY�6x�i���+�S]�&п�̧6��D	/*BPL�d��h��O'��5 [8Q��Q�%!���3ݔ^�1�*ؽaZ���y�f��*�;��S��̆)��Ʈ���@&�bA0`���%{��&eiiR�����v���?(vթ�P����G������K�p���z'���� ���]V�i���˯&ON��wW�g����8�y'��1���2����G�K{I6��'�M2(��C�Ej�#;�wVq��1�]'�<Ѝgޑ���O��o����_eJV*�hxل w�y5�6�[�j>�����c�L}�]I
�@�#�Ĵ�noi8_��Ad>/F��Ew)�K�1�+ԑ`uSW��'��1\5K��h�t3�@�#�&����iߛ�x
���^����;ԓ��������O��G�B��yvP>q���ֻ�M�����1`��z�tr�
��� �/\��2'�_Dw%�@ )|e�O���>����e�f5��28���LY��Y }���a�2�[��r��O\ʙ�*buQ�����	� #vL��[ 0pv<O�o�\.^5��J�"����� O}����v螂n�jj��zPMSO,��_t@s�4����<gGe:��'j�+O����M:ӎ�F	�zܖ���L�5y�{����C�Ӄ����<Cd;��&����v��RL����)��чw�����?r�l�g��3�	J���&��VfQ��o���*�r�����2֠���{7#{C��o���;�C$eN{����q��E{�7c�4�eo���"]yU����F��\��G!���̊�Ć�#���|��NFu�p�F`�>��hl�lɚ��@Fà�ñ�'rں���+T!�ϛ��w����ُi7=ȇ��A ���տ�Mޕ,�����A��D�X�m����}��4z��(�W�i��*�Lo\�"�B�x� )2d��Ĉ�UNI�D��#��MJ܅R5��(��+1�q2��8c���	�"�K�4�o��Jk��ut}�O��h���䆆�fN=��qIt��������9�6D����A���)�l�ެm�f�Qi�(�.�,�TX�/��{.�0t���N��<|�
��jw��DoH7�*5E3��K��W��Gsl��/B�oF�� ����E���~u���}%3��� k��4n�'Yp*�5�p�ݧ�x����F��I���%� bS���Y��f�!q����{�*�|�dzT���[ȎE���̢�wM�$dpB<K��g�S/H���ƺnƻ2��t�;��LBC[��"^���01 ��d@�PZK	r�$ K�j:n�7͟�)'��Jr�z
d���F�DNz�8����lDkN�@�-ZR4xmg'q��q��+'�U��ѐ%��2��@�-=�T�n�K
a�K8ґ񅝣I���n.��򥓵WT�)IXo����k�����-��9��qq���sp�*�C^��s���g�G�D6�ϴ�Ց��3��;!�cL)���eBb}�׳0���嫂��ָ�.�_oPZ:V޸���M�F�7.1jzğ���A��ˊ�"����ҕw�(5ky����W%��'�~�ݦ����3��!#f���t:T��	�n��RE#��Md�酾D��~�)���8T��zX�K.+i��iS����]�\�4�ŨA�^�2{S�w�kb����V]7"�~鿿rf`w<_0L�hTܯ�iIYb��..��0��C�OZ^#��{Ɣ
��Hm��,��2���=$���_f��q`xP��5-�d�eW\u�8ř����ȳ�O��7�����a5AcM
��3m}Y���
7k��.I��$ގ��:`�)��ElJ[�wDB%��'u�᧗��'e�� t���n�	J@�$-�����m-ӊ,�������U�A�;򴀧_��|�A�p4p)�%�X��n���Q�n���ĩ�Y��W�1�?��=�ou�`P�Q�K/eD��H.��#y��s��������n\�ӧ%��F4.�)+�?�03}L�241�'z�d�C/�H"	�͎.XZ�������٧�RY�ޱ���¨��ם�v0ѭG|����+X���%�;B\��`�k��
��&h������e֤���@�#x��j7��6���?$c��^���(vx�t�����_�A-���.�!K  R�++7UQ���AϕL�oW3R�G�����΋CN]�*}�/QW��҆�;�ު6���(D�+�C������;`R��E�Ebpf}הm��d�I�8�⿌r��g-�����ݧ|���8�{����H$�������_��G��"�N�M1Zuˇ�H=�
I��'�?�H�wk���mz�V������;����K|���M����[�D0�ު�AmK�-�r��E:ϑ�z	�9�<R�ڪ]� �}����
iǲ�tyG%2;Ąv/]y%��cf���'��ퟓʹ�O��g-:eg��w��ޏ�c�d�$���`��u���,��QaT
1:Īl��Jx�F�-[����Ց�6J)ZV�Cy5�^]���Y���>6`��ɚ�b�E'!�[�.]QM!�:д�{B�C���`�T���7%K�2	eMG٧���m���������@:v�-�L�忖��(U�U�����/3iv�m��k,��@�)�#d�h7� ���#�s���Sڟ���)�˯�E/���MWC4���p�C�Yq;����U�\8��`j}����'��������ĤI';ky�%�������VM�#'��2b7������\�W�K,3%k��^(����1�t$4=;9&kQ~����&�zYZ���W��~�1�>	��J�t�O�]��P%�$R�#����ju`��˂6�2{���&�����cT���Z�x�x�:i�3�q�#���Q������Q�����<�p�:���}33@|�Fs2�Q��E`�/_(��$X}ڄTЖ�*�?�2w/ӽ"s����J�W\����ݚQ0�?ǋ/7�Y(cj���AW����Yh�ѭ}_&�i�Q9<�~Jx=(�[V���5q����씏>
�X4�iD?jQ�43(�?/��K'33o��"/j�ױM�����C~0�l��v^�����\53D�"�9�%Y{a���B�j�`�2��6���S��uqx�B�,��d��T5��>��
%�neb����^����M7?I
_����i]�$IFc���xDt� ;E��aYL�{��W��@�𦒵�ؠ�5���=i�<<�>�8�b#���t&�(�C�x��,B\�5E�c��t����A)T�(^�]�Xǈ;|��Ƶ��y
&��
&M����ST_Al� �!.�8���ӢrP�p�8��Mg�d��1|�a�!P4���ì`��5���U����޴����*M��	��F�|�w]|�iS��J��o.{\RQ;�i0\q�Z�$u�����@/J�݂-xC��9��QW�K_���B��fn/��?��`�]1�B&Ec����I���ƈ��0X�%��>�&H���M]#왻��P���(�W�Д��B�=��d��% o�WuW�|�_�&���iC�01�=���+��"�� ���/IJ4B��c(:��w���>tOY�Q�:��ۢU�r�q�fg�=�X:�"�n�Ɋy�u��nw�{NG즻�3H�L*�}t�b���{E��R�E n�4g*����ʜxJҊ��b�����	HѾ�#q\Ϝ��r���ڲm�e�4�e���(+	�QWQ�^��y7͙�)�z���
G�j���;zq�m=JAT��/cC�T�N0��%� �=��P)��S�w��d76�Z)H��؎
��h�:�������S>su��?B?�I����D�;��Ω`,C<�#,>!Ín�&�Z�2!�y<p���,�É��x)��U������9�e��Bã���,��,q�"�[�s��	Y(�=�����k�'��Z+�<�d&��9��[�m��O���}	�2��3�E�Ͷkؒ�T�f� F!����a[F�[������Mq
E*���Nbw�)@�D����X�E;�����k��ViMЛ�BHO&�Kل��~�1�p[��1�v2�Q"��k-��?֥�ϻ�E���c>8}?���o�xqf�u {������~v��;�A����J�^G�C���c"�rPU�M��a��F5�/Xs��)+6���M��߉��I�~���%�.yH�0fF���M���3BߛJy���M�xu�`���}�C�Z	��s�Ռ��WrQp�V،#�ɷ5�,�^��h*u�d��	]̧�� ��E2����ɌO�/�g���V��`��Z��&݈}hV��,�mN�Ї�6آlVse�"ע�I���AD��z�Q���+fl�ڒ@�H�8�+[�j�~#Vy�K���%�K���#��e-P�'lpW� �dU��.�*��|�:�{�-5�L6�K?.J�:�FW8'ؐ��Q.�w��՜��eMpd7W�+Ȣ��g� _$a��&����f��#�l7�X�KIܳ�y����<|�\�S�Q�붡��$Y�9�!Zp����� OV��L���n:�mA��G�$,mx�W�f�)'��/�T��.O;�9�J(�}FL*b7�[C���;�-�@Ƨ�
�:4�\��A���1�6�#�r�l\_�c�T�V�C/�\&�XHP$ח�������d��k�Է�����;yqpF�!-N�"+*{Y��� ѣ���'��r�?��ã��J|j�kR�uG���)ҵ�`	zU�o�s��|�?ea{����$Y9��9��5��Of&\�{�u�|n�7���F-,�H���Nj��=�S���b���,���R�b� B+�.�C$9���%������c5ˠn�5�{��_��<|vp� Mb�uG�Q=-�L4��/��� b��)-�!r	�|d�<,6i�:ې�c !e)�+�� ��@{6�YY��9�����|�A'*�>P��v_I����N��m��� ������g`�I3w/�!�6ck%�go�%E{M'�*�N�/A�Ȯ	�1�_����l0�W�MoV1n\�阘�Z.1r�d�`y��[ł�DT?s�"�.m���.6S�71���& Z����2fK�]V�wp�~,�&����[�h8����~�2R�^�cp�ƚ��@U��R��D�clb��Q�G&��p� 2�$�Qk~o�+�?i��[��5N�w�W��NH���ı�ρ�[_��WՔ �-��h^�土W;�H�ro�z* ��!��\��̨�#ES�v��h�_[$N*��P�D�3�����C+O@U��.%f>{���$��d��k�Wۋ���~�WJe� ��������X��PmZ&s���
���~x�K6��Udy������(���5�V��<�ކ��:�|��=}zH߽�� �f��؇�)[��Jy����fA�Wg	)r��)�7�G��УHj��!n�"��q��1��\�g���g���(�]�AQ��k��ٽ<���+��4�Am��-T�gM��?��'�q������;��Ҵ����i6h&1ʇ�X���Ŏ��|��!���(�-Ӡ$1��UD�b��U���P�t�Cq�ӂ(Gz9!���h�u�ÒjȠ^%-ռ���-�)R6p�e�Z*gL��I�,��L ٴhD{<Zp�ꤼ1�� ������ϻ��s����gcw~��?���qH����ݞO)q�ʵ��E���t�p��D�_i��γ+%b��R����2�YҾ��O�
(���O�d��VB�ڴ:����.B�1�B�'x��+��`������-�\�^�Xr^�b#�K1����[�-�k�!��:�JS&C�c��K/�Z���of��Ny�c(��J�8�:5����e� �X�k@�+5�.xn����Ѵ(���A4S�ń�0�eC����
�g��mM�k Ϭ��P�9O���0⣺�M�
�E΅��{��������X5�,0}��?Ps���Vr�Ѫ����B�J�#)��%{����� V[��������緆��a��ݍP#��<eV�zW���-rax]�?���qOLضb&AO8>�P,Z��:�K{v���F2�E[�t��{�]F�ƅ��h(����,�o/�I�������[o"���f^���=�*JR����ǬC���u����q$�	 �����V]�g�C،�A�%vO���s��2�VԐ˃/�r��S���7U1��XoUOR��\8�Y�	_XoQ#����Nu�v'��-w���S:��2�0��uZ�7�;fH�.W���8Q�h	��	����LR���Eg(���?^�dޏJ���-O��(�!}L�A�mH�ilt~ջ�N0_}�y�����D�U?�k�;�^y����}TЯ���\�ٔ,��8#2��n��6gsoL�*�(]�x4����y�َg�c%�К���YM��i1V�ެ�1�NȌ�]�2��pgeZk)"b[1\j�dQ��=1ߩ_���"�8�B�e����"�}��[�#+�d����]���X"�qI=�.z}f5�M�Һ�AlսL̞���=����p� J׾ בzfa�����|8:�&.)������y�oy�/cK�C���?�3(�K�����Ӱ������ř=0.��B�Cpa�n�u3Αs�H,��y*��n����z��Iq˥�H���R6�z�*!_�e����^y���r
R"�/�����T�O�(r&��
�Ti�J�Gj��Ъ�D�����O�
����Ҷ[ϱjvT_�p��Qۀ�p�t����x~A/0���L���B�lc�{+(��ϩ����m'r��A"�5�q��nK��zb����9[��>,I�v\+�@l��b���L�_h���Σo��4*�7��NIU�̲AXU�1�˫
ٛZNai��ƶ� T���/��Z�H�<�ҹJ,
Q.@��)i�b@r�bRN�w?c�keパ�C �GzJ���h��μ��4�f�(�}|ȯ���2��ݩ�YQ�ve��eW"Q!�F���4��R�y�2<�1��??�� L̒�?C�%y�Pc\743�sc'��e��gM���P���:C�������j�Չo���#�n��R�v�����Ze�̵_F�槇!��j!��W\���6����z���.�������&����.�QknX\,�$j�˺�q_��4�L.�_�IU��#��@�1��7�e��=z�a�;��QD�c��$����(g���<��:h�I�� ;RYuF�e�o�%�6~��7ٮ��WVN�:R���[���%��{OK�S��V6R��*Z"6��d�@���p�}��`~谅�����R�ht!׺�z^�N,n7^x<:���c�/: Jы����cs+hĩӐYS'�`������P�"�P���+SuC�b�k ��߄� �����9"��sU� UQ"񊕮��>"���rZ��y��}�$ �JT����x�/�k��9Ëcm4���У�W䒅$�ohZ�!��X�� 7�?G@e��qk?�������2mM�C�#�C��H�<�1��+�b�uL=�VA\=�=�6u\���gZ?�χ�i����*u�0��/��Ul��s���1)n}*f�$�|�c#v����Ǥm�vX���mG����"ꢳ�{��{��Djla��A�6�w�&G@���<�eg`\x+c'ۊqRqs>F��]7�pR�>��d,�
���sk��Tݼ����9��i�'=��I���Յ�H便�5�FT�3a�u�7LV��Nk�0�ȝ�Li����Ř1ݥ{K��?T�1+�	I����Wȁ���N	������
Br�Y&��sS�;�����B37V����94��C2}����A�KV���ɱ;��š����[��=���z��4*�ADe�Rd�/yJa�w+Ç����톡l�O>M���~�+���[ʁL&��ǰc<|�hZ;�r� ���a�+��F��8���Nh�L�9���ʲ�~�i��C�3)k��=��Y7�������e)��h�*��l��zQ�\7�,����䁂�(�t��D|��mC3�ڿ��gΊ~����h<�.�0P�n����$7]��#�v�l��
3��[c�D��' o5n�ç��顎�}�zm39�D�9H�ʵ�o�#���\�-�`��":�Crmy�<�H�p���oǂ�k�=�!�<��ǆXs�j̓��AZ�Z˒�q���"$�9힆
�rπ��u툫�ײY %=:�jm����ۇ���.G�jj��?�:�KYK�A>�(��'�fV�V9'��A�.}?����L���1�,��J;݇�N(#�9d�e�u�i��!��fJ��U�����s+؆z��@��!�5���y/������$�|n(�9�$\i�c��Sj?!\�w��rj��7�_�f�{I8&e*�D�Q�\A��) :~����P��$7}`���ڥ�������m�?$�[3���4�=�@�5��J�!����ˠ��vA��t�c�f���k�X���o�)}����r�Z�1ߝI�����P��"�Yʣz�!����7�=ʟ��i���:�[w�l�2nW�1f3̶TS����]�'J��s�]%I03�W}΂�(�P��ؚ���;��v����/�#Y�\:9Q9h�ՄaWeV���lv�*"R�e�`{��"r��7�7���J���$�ܪk2�����x���av���w{I����]����+��Ω(�*���i��Ո�~룞9Qg��0}�T� ��ɭe�+�����l�]��s�d���� ob�uR�j���ч9������*�gţ7z��'�5/)�C��z��J�R��e�Y99�U�|����G�H�M�]�V0�	q�xiDKq�oP)2����hZ�U%�2@!�_]�-��"e��,�H�v!����f��P��l%�ݤJH)#O�Y$=RS�[qB�
����z��Ёo�'5�_��&^A�w-�ΐ<�������;�M��\��5�٥����oTah���\�_�0"�4g�'��AW�*�1R\9����Ъ]��c����!�F�G�/%���K�h�EXD��
2��:X������c	�Z�<� ����EW]���E0�#q��vCY�K��kOL��Mҫ�1�\��pҶ{b�J�tV�A�>����~+<�˄˕ft�-N�w��( �N"M~��}�v��oHf/��-n'v���V�S�*�3�f�&��0J,���ˌd��w�i8��5ރ0n Y�B^6�� EF��!�+�>�fT,�^M]�����_6
��9wb��4��}D�;�Z6���}R��>��r����=�!d_� �w���o줬fУ:BVC�v��!(�R7�!�a܀�Q:p��>,�MO������Ҕrrъ�o���|Su��|u*^J!$HMX���(��W�~�'�ܒ��y_F�kgn-�%� �pOM���	*�`�S�M�I�\ ��V�w���s��&圞����5�W�,`sf��>��԰=%��z��X�L��/ [kE��'�w��i�J�UZ$í[�&��Hs�������,�A��/���{�E���G�y��G.E�Nq��<��y�݆�Ys	��7�)�A�)Y���4X��u&Ǖ�]����4�7�d+�Iw����Ž�X�ͦ�ol��z��A�U��㹝U�(٬K�A��<z�r[�<���>�T��L�a7��	3����b��jr�>�3c�UU���v�2ץ�Y��r��g�| RYma!d��N]z�]��R��O^%q��<U[;��k� �=�Ƥʪ��g�tyu���M�z\0˯�s:�3�0T^��O��p6�`l��W�/�N<.gΕS�pK�ҫ������������%j��
L��I�+�8�)�ۘ���>�fj(�@�G�$h�z2TB�xsW�KrɘxtH�i*>'���������A��T ����u�W6s��,x�+�C�W!<�%�]d.�qN�O�B8ȣ`�4JN��/l��L��?�d��x��	�1���=v �13�a�?�Ե��$F�S����������u�#g�M#��'zq��ݿ�������wO�*xz!�z� ��(�̀"l�-�D���-�U����%TK)W�~WU�^�@��ߞ���H�О����$�5H߮pDy����"��=�*Ҙ��Z)מ,$�4��F10�} �*�������� Y����P�M�A]���x)�� ��s������^��V�ak��|zLS�j�=�еf��A]�I��l;�эG��R�&�UՍ����2���zx��>��DR��~�� #A0��Q��q	�i�B	�@��r���v7Dy��N�!�W"��S ��ܷ��;F�=�;8��XT���<�D��)�j�xsw�\���ҋD�Zjθ��b�!"(/�@��[b.��xuo%yi���Dg�� >@���D��IZ���D�l��Sv�Qe�%uX�蔝��q��9�_�/���� &1:�.N�P鞕ؒ�jE�Ґd��튌

V���k�L��������F3]����YA��J�\,��p�R~�eErۖ��?��*�{Hڮ-�ٮ�����u�����_i�~��;��ϥLyˬ������|wL�n{��F�КØfSKh��@�����O6�C�m��'LkH�1�M���I:���At��@�L$�c����A �ρ=/Q� �O���eH?K�T2KM�~��2@$�/E�d�u�~�۾�^":��|����J"a\qY���-�4�xv��乱�
sA^R��)d��=�C���s��9��r66u�jQ��Jt���J/վ��sdzղ�������yV�C�ܧn��E�����s���D	������z�Q���NX�ڦ���}�	��zȸo�?�`�%>��;�V"c��%d
�]�7�%�?u?�9�R�l�>c���Y!2.��}?�?�9N��R��!C�u��.��x�te�������dB�ТXzp�IP�- ϕp��!a"*R����[�5�O7F��xin4{6�_�(X������9c췎� x�z��C)6���\˓2@I���x�<�"��,�	t*G�Sbz���~������f�/Y�<���A�7�y��D�)ж%ul�ߐ6, >�}1� ��q���6���5�ϵ���������Kwn+�%E�j�0_����&��7�|)����<0޷�������h�o��.m�LSb��G��|G�ꀐӎ���j�Z��"��ЪT&����������5�A7�Ÿ�����ښ	�]Ù4Z,�q��m�}7yf�E��c�(rd�pCm=���1�7��*����{��z%��A�5g��_*h5�lr}�o
!:h��I��(���LSLFA��p��s�iz�@%���n���6�O���ؾ�L�Iy��w����#\������k�z��CR�Y�z��Z�!�p@��>�Af�>Nϐ���Ip,)� & LG�M��}�GH�|��?�0���o��w�B�e�
i��ek	��- �Ѹ�1E�wר9R˶l5H^�^�/aY]� �"���szׇ�9wړ���% kN��D5�s���k�Y����ƥO�]�=K!Ƣ�y�E�6W�6�O�� ����������m��d��h�2����׹�����Wpw(0)�zQ&�vU��¢s�e�ˌ5ޭ�6�޿]�GO��q�鑡��t�,��B+N�d���5�upNz�Kj}4i�8]E��V������ƃ�y�4�44IǰhB�}:Y�����QﮆTع&Il;�[O�*���}���o��̚��&D����O�� t,��^�P+9�B��w%� �hQu:�F1y��g���֪N�թ	*����_Z�!�qp�d|��a��/-b$;w���:3I�M����j�㚙�P`[�>�Y*F!g�vn���^��(ꓛ������-չ[E���Ay������B��*�n�'J������]��w���I@%+2� ��׭\N�i���k��҆���?�}��e�frIQ��B�J�ꬅ+��㟋_�E�(dJƞ��ᦻ��dPJ��"d�%S7�V7��'��3�q\���Rn_�{�����{����P���r~&�O�%Zq��P�]*���<��|1ө9b̐b�A�Gf̼��şSl[ig���)��#
��4�[[��<�"���t���=�J\��@s��}f�ذ�n^�:��^x��2��m�W��z6����[	<�9�*�Qe(#$��Fųbt�����2�6�{���%������o����>��V�Ȇ9?}19~�n���Ā�~��+~�â�ޣ
Y��DE�A[��@\���1׆"�G0x��ӧZ�	���̰�W0���N�݉�'O�⑑8�1���$��V���p]+�M#<�K�k�N�tK���w�
�ӡ*B>���*u~as�s�z�HFF���"�`���qclԳ!b ]��K�O��dН;E���[��CQ�6�4Fa�>B��āTw�P�*�$�g-�l�c��2������3fȅx��9��?n҆bZ|��5\�~g�В���(�:1�w.c��܀�������/�H��͘�x`�=֢�Ŧ%��3�?����g?�3̉L�0֤�[9��T�r�_ŚTU��A�w?"�����L��_�1��j�=x���l�=�+V��6H���D��@׏Ԟ�W6�$�s���q�*���2@�l�#Wn�<ۆn|(;Wbj��ǺQ1��p���8hcƺ�����B�-�E%�-��>��Rx� CSs����ײD�r�C�n���OQ^�/�J����y��ǔ(sv`�l�������
�WC7I��ƍ%����M�U�v)� ���*��Ζ���b�'�;4����SW�r�%�ő8���"�bT~��኶A�S㛿z�:i�|$�K6)b�]L8V	W�@��x:(�Ԋ�Z���ǔ�G8�U�lTOmG�i�-�'��H_ϐ���P����/�:Ҕ�c�V}��G��d#� sZ�p-����L��Z`V�����[��H���b�C��}}�b^az)v�eay~�w�s:�˜3vF԰S�?��&w<�o&�<�\��0@F�����}���JbT.�k����,֚抄��|a�����B����1��҄Ai�fCk���-��%��?{�������W9�[��s(f�480R�I����a��<��좍Ţ}q�5����n�R�V�4\�p�	��0$�m	��IW�� |5�l:����t曰�#����J)G�ϥ�F,t��l6�8U��)�]��M��!<c8*�/�
���;��gS���q'��F7gK{?k=�atڌ?�<�j�{��+�紐E��y8�3�V�I���V���sHj���X��D�8�J�l�j��O3&^L֭��~��O��Dj���t '���+��>��K�_>�]��l���@�a�}����\�1��9����/�Gn�Djc���,-�N
ה���Eq��o{ ���R6���i�SO� �)�~}L��ۦ�|!d���d�CO|����ׄ"� �Pp�Mh��n:]@Yj|<5�v��������Q�ŗO�Lb��ӑ�����QQ���|�~� sY�1����i��X��`�	���uҏ�;��?)I��/��K��qWZ$�y�wZxe���M�䦧�]lқ{4�넒��Y1��݇ a5&B��8���djyo�FKxlV�M��ݲĴuYE���Y�i���_4}1љ�ȸ��]H=J>�/x�T��u�}�ߏ��V�����Х�n]4���u�vJ"���� !������J9Ƈ��dX��J�w��d�xp����,cAwf�^���6N6�m\�Z/sR�	�Q�\�圞�g#iĀ�Y�I��9k[}��?�%������c�璖���A����X���nB��r��ET��� �ڒ ���ڰk��Z;σ�U-)��#��d��&<A&�F������V���#kk����
�08��%���S�a� _-���7�#A��񤭼उk$����ر�Ss�<詜5���'9+���G�z�L��<v�����丒xڻ��L}�SV9�k�,/Y޶�Y	y�����~e�Lw9�w؟+��`g��V�P�@;n4���q�w-�Q�fZ�s�������+\}�r5�c�SG�hJ^�J�=���x�h��`�$������2�����a� ��	��1�t�/^�46��Y+��,�KB��Z$��Q	��q��oR4�=o?p�\N��J����&�[c����AOnP�4�f�.[�i��y"�n��~����XT���HZ�T�Z,i�'8��}'���J�Eɚ:^�����-#��������W��Ŕ�L&̈́�8�*�/z�<����	'+��R�Xƣ������;��Q�?�`:^}�@_m�+��T�t�;�{��Am�H1���W.� u�n�E2W�np�s��Ao��ӡ�"	L�md$�<�\���G1�1����3�f%b�4��Eܓ�=��Y?���M�y�Yo6PVWQ�仙��s��X�r5ES��
l|�`��{ڙ�L&c�|V����x�9����IUm�j���HM�TǬ���(�GB�{��C665<��[�U��;��/U1M�o$�`\u�Rό��ㇸ�vX��_L��Y�9����l'~�G��^����B<kd���Z�ET���T�6
���[�=�������X�6� �,|�@9������UBs�ʒa�;�YX�v��{�4�	iB�,��@e*�����eT*'��t2��i�3ʁ5���$L7]��l�y�����Oߋ��;A�%�K7FRP9i�\"d۸ �4�Ge
&��o�����Y`���9x�^�w�E���_n�F��=�rZv+�3{&4<:����3��Dψ��g�_d ��7��8%L}�7�@�y��e�e7��p�'�Ҽ�K�Q[��ˍ��b��ͽ�-�9��+\<7V�)�1�_,,���~[��\}� � Zs�<�+�xt�Ba^ ��A^{o8��Ӆ��-_]����J'11� Ŵs�+�+�{/��("�p�A��pI����%�[,�`�����^2��ׄK+����s�;��`E�ׇ�4ΛR���}��t�$9��xRS%whF���_���J̬4�����5T��ԇ�=�W�U���lh����%FG�Q~�
�U�#Mz ��XXC���3���^K�9�{�;&�v*0{*�,�(�E�0Z����� P?�F󚐪|�t�E�vma�N�7.���v�����렋N�!\f�����ZG��h7}��1��Q;@~�lfM e�=�6�Y�V���uK���eʻ΅������u�ѱ\�g�2�ӏ��W�lG=W�h'��̖Ă�^Νq�^��+��@ń��P�}j�( SbKx����S��o��v惷��k0̘Y��L�� �6�v>�6!#^�g��K���{��Ð>�%�d��C�}/Do��KG���t�6�"YCȻ��ц��A�|�3�������V�C�=jY ^F���l�k#������Rr��	�kI4SK�}񷑧�Fr��\���f���@�X��(�<ǍI��;G��0�L�-���O\
�	8�4z�=,��λ���u�qr��`^��`���?�򽂙�KG�[�m��<�B9O�[5��>�/�& �>����=W����>����V���!���Gŋ�#���uH_��C4�D�.��ѣI6#�#1�H��=@�_b��j;/�(�&�p�Wm;@���C�#�8�����#��'��uJ���b('�_K�k�Rު-k��!<�u�7�܃��WL�+Q�m�-�Fa���'�{���tț(�
���y�*�ho<e���Q�$[@"ܓ�0��56 krg-)���i�����JN�"�j9�XK�:�W �(C�u�v+)Ѝ�)�q+O��_X��o�z��K�h�`V�3�yL`*@���+�Iln�(CݢA��Ц��U�!��<!�����<3��kk�~%�>jS��^�Xc��J�ĆNDd#��]%s| ��ʌ����|�5�^�����a�� fS��`�2"�y1^��WW�hm�ƙL�%���i��dvβR���]V�E��w��X3�ܻ2��Pd����M�������������H%�#�m���?�~+_��"�lO\{v�k@�_/8b������!���C�1��ًl}k`X�\Ф
�U�!�"�����K&�n����X�fy�1�:5�F�,a��5!�\��0�U���g<�F%H�
����iO}>���g>~y�=��Ê������ͅ�$��h�m`���
�ʥ�hc���?��5�4n�Nא�-H���4��1�$֛^g.�Ł��۬���{w��B�+#�}�42C��/�Ƒ��P%((I���'%�t��[񌂰�H����q�ߺ��i���ƹv̒���`��x �����Ø�'��)���h�J��v���&ɇXx��׊�����^�_MX�2�1��z�e������r�o�s��8y��V��/�Wt��ęaX�Fb^9�P@�Y�-~KK?�+_W�2p�r
�0�*�a,9�Nn)X֝��p~%� 1U�i"��fʓEc�z�i��Sb��g0}�8���mNʴЩA�c��Dچ
/�_�J�c]�����0�6�ᵾe�i/P�����$Xƴ���|~"$���IWk��ɬ�-Oq��x�6c�bv���C4�n��iǄL��/K�f9�C4'dI����!A�j��T����0��`��}��/����>���Lx���c�ر�I�y�!�M�Uϫ|
Iy�{���"J�;s(���_@���ȧ��}������o���Ѥ�^oQ;��, >�K ��7�tl�J\���������d��N)�窽Bܗ�@;hCK�!3�@�Κ�������{$��x����&7�V���٧p���j��	��'�_��!����EJ�;���AE��o�����oL��� d����8&�/�9�^^�'~���xw���W�m���g|�C��g�N}b,�{�^�:��<��V�F�!�����/ͪ��.��˿'�Z��s�r�:����pe��ה��C[r�z刾
ϴvi�� f��^���d�ZR�	!�� ]�F}�0�+��,�!�]D���X)6��y�kW���ֵT�/GR�gTJoI<A���M�0��bi#
�������/}�Vʱ�u�M�N��f��[,ZWR���TS/��C�� �\K�����ҡP�����PT��
Ƀ������+�j���(W"<�	H���f�~���j�2\������e
a`&!R���zy1h3��{)ms�4�`�O Ӆ͙ɱ��p�o�ra�#��28wC��Z��f��՛~�I]u�dЊ
x�q�x���O،mu�?�b�|?�:��UG��ĺ�mh�-�G^�a���=Lc�Ę�g
�A[����bxڌ��/�\���=��(G�W��!L!7�ۄ%����?��+ݥ��%Ț���Ұ�]�P\/��dIT{+���ku�$��C��N����I6�MR�
vӀW�l�XF�Z��}�N_�-|-��J����6(����	��^P�%��A�Bd#O �7E�C!Ra��U �nT*��4�#v�Z�Y�\x�E�Ԓ�&�����F�x�<��Jx�H<и�����3v�>Z��Pe�Iq��n��Gp�7B�=�a�şB���F���b���ݙ-fߗX�_�uiѱ���W�w�+~�#4�L�sj�P<�� o9�����@eڄ`Gܼ�A�c�A:��12�->N�xm�y�=�x�M�"��� ¬���"�r��$�����A�vlC9�|^�Fu�d�Y��u�mt;l�ܧ�I^�Ϋ. �P_�kl|��;�1��V.3c�\者���9%�8L*���XL�R�^^�gR��^�6fj�7��?�'X��9�Z" >`�3l�'ԩ�U������N�}7�d�1����@ٹ��vg����ѳk��h{�]���|��c���. b��G���ﾅ��G�F0X��#�
𛯠h8��ꝃMB(�Vr�z{�}'����2��!���~W��5ji�}y��b,�y���j��/����/N�z��x'>�Z�������0�H��s���'\�O.pz�,.��0���?0�=�kq���#������8i^���kV�S���cC�\/�ћפ�������2B״c|D08�X��m���G���BUo�H��f��h���,����R�ť���M����
GP�]�S@��׽�j����r^6D�R=�`;�l�Ղ�Lo� ����f�Z�e�5��b 4q����LV��V�^"VS�8�6��k�
*.4�^�RbZ6Q_�Ot*�q޷8�� Y�:y�$�#��E�Zl�ܺj�W�ц���y Ė�R
���w��R�߂���	�Pa-��
^|1���,�Pȏ��({�V�"o��5O*.��*���@܅�V���5>��wJl'�V�n��8�G��q�x�J�F���>V�]�LٳM�WLvԬ��*���\��Լ98�F����Oڔ|h]<'R�R"�QR'5c��h3�f��&�*8��tU9�#��z �}�I�$6
\���?���\p&�/Do����A��L��o7L�>��/q@�M�&�d���ջ��N�i��0g�.#0���P@�vf9����SEx��_�.<��(G{�[��P�������Gu��Rݰ�J��L������3d��bW�R����x���y��L�0F<��v���5/���4��4B���B�w�Ph�iX�=�G>�*mY����*Ip�Ğ�оqT�<Nf�0h;���(�b�6��L�kkz����T��z����7Mt�|�#+7iM9���~�W�O�]9@�&${d��o�a+���ó��"ɓ�D1]|!���*1H����z2@oW�gI飏U9��g��-�h��h�VV~ދ��τ���O�-U���I�	m������3�P�4Y�J%�}b��Q����!8hT.����BaƊژ�qu���b���͗��3i�6��%園$�����FrÏ?9@;'��B$����GsJ��;_�m$���HR�Mɭuڪ�wf$
ez+�x�U��G�Jh�׏�����y .��I��.��h��qRh�<��?�)��7����z��C�\��D���M��K�l��}��9�p��DP�=��$&���$����eg �3�[w�� ѕ$;�����l~kB� ��ʹ�4+P�1;���)O�'��f�Ԕ�̽��{p����8�5��U�D�s�mt�|����F����!?o*qv���� �WE���i�=ń��rr��G�# ���p�k�h��qI���"˥����b�=��#��C��E�"���z�#>po(ˎr˔y�j�'�����a�g�����Lw�C���MO6���RD���?�h�m.k5{�#$Ҳ�NFò�[��2j�.��q�� �+#�\~�����$��
��ۥ�(*���!�RP�h��.���m�<̃�B���'�S�'�W�ZR����8�.
m��Z�tHKp�m�2dɮn,O�u�Ȇ2 d�������v	��Q����`�-�$�sG%/$�4�f����ϼ��(��&���!�R����j��82M��R�Ez��MI����TV[\�^����S[5��S�0�-�61^{��{/��_�7YŮ��6fY�a3}`=W'���Ԧ���M`VX�J��mF���>������Z�62�UBg۳���z(f����� ����*d�`8��RA�X� �2$7���*�o˂�t4��Z����Sa���0�@�,���h*4G���vtto��9�� LF�'$84�M��}�2O�e��}����.�v�PL�y���p��90��6�F#w����E��ȓ��c�T������
�g�M�3L]����w�ODBg��vh���iM�.X�U�8�8	�ɬ��|������y��b(��sZ[1Z@�d��C�<���G�7_ج^�t��"!��v�(cЧ;YBz�UZ���q^����-�UQ�:i��{�_UV�JV�� �6C�t��|����o��Z7 �M-]"�̅�	�<_�J�[�޾�%���%W���84"�{�̐�vJ��KJ�-��	#��F@,�V9v�1�O��e�H�TΊQ���"��℈Ĵ�� �����Tr�N|�}��cTX���V7}���<'-;�*������,5pf��Rf��Sf���[� B��AI^sl�>U�?�Ұ���j�{��UZ�8�?�Ho=����&I�!��T�~�2���aN�Ǧ+-�z��žD�<U��Ѝ3f�yN%Q���}WL�g���%�� �3��BW����/?P��y��1?�K�����R�mJ
1�u��b6�fFj'<�g�(�3�����Z�n��Li4n�,l0H�\�i��L�;[9�19�i��_ǁ��' �b����F�j��Z�c���3�\�,�0Ó�����6���pj�Ms�8�D�=�k�;TTmc����(�F8-e5�p�0���k��JO�`nϸsF}�|4�2�]3��]\TZ"����j�~�\���M���k'�Ђ~�[�ȖA�PsĊrq�"�GS� {0�����Vii6Eu��ϟ� b���U$y���a��5��KW�x-eY!�� �b���Lxa"3�����,�X���Jvr�tG�\��P2��5͠�S����l�;�k���Ka(ɚ�g9�����Q�f�QR�VX��G��G[��Z���$�˶b�$u����N�ZL� �ź|P�갬�w�f���>m�!F��{�$pu��y�����/�P��k�W"MS��+r��JS�N��ћf�Y�B}�~J�a����k�"t�'^[�!��,��)h��-�^p/�uT|��G�Pu"5�
 DG��Tr�5�5�1�(���82x�t�(�I�(j������Տ ��ϭR"X��d��$ɋ
���1@i��w�A�,\9� ���̯G�Rڈ�/�E��ᗊ�9�� \�[PDO ��OŞ�]���ho�{�$��NG�<��A#CmF�������!)N?�"�b�HӸ���<�C�斄����]�B��k��.��s�?�)u+���,�'N�=hA�B�M`�oϡP�-I}�~�̵9=ؽ4�v�����ɀm26�-Y$-	�Di(�Ş���1���f��(�-�8��z{/�3DV�Ƽ�����bv+�/��_ŕ������g)L	ˈ�dLE��̊!��)SN%k�]>�����ϜJRO�g*%���ƹ4i�����!"o�F(c
��E�1n)�+�C�����)�e}yHEz���v�3T��]�2[��v+]�XY8]���UN��K_e���m	�����Ziwd)�GE55փP�Y\4]ǡ�~��
�~P�45d���=H6�	�j��#�Aq0h7Q��-��${�*�Y[z��r"�.$��袬�e���Ց���5xC�;qE2,(q�,d"4�X�nD�f'����vW��W��9�H,��jg:�������틺������<1���9�܏H2�B��c�E8X��R�,�L�ҩ`���]^��a�
�lug$� ��V�Ζ�㧉h&�ㆵ-��L>�����`	AL;�^���y߷N�K�˔F��{7�����Ѯ�:�Y���?����<\M�\�f��fP�ܷ@�u�"H��5�'B8�3Jc�|��m�RN�A��UO�qu.�lըULE_
����j��]#���ޝq��������=QL�*"�`��Ùz��9Tb,#��m��l�TU�0O��T@���qK�;E.�.��r~��?_���'���O�,�/��N�T��o��^�O��9�p�:׮�e�0h@�P��9� D�˂��/_5�3*ȗz�='j �4�N5,t]( 9/
�3�g�� �#f����dκ��Egm�4��̸��☇����Ug:���k�I��*y��p�6ݾک��Fy��U�	��$S ��N�(M��2����8F8L=�+���YiA(��Ɓ}%|0�B�0Q��l]��#��}w�`�i�����!HȦo�]}oF���C����$��УD+�OYn���7E��Y�[�3[�� a��>򞋎`99�)�B�S�/��bL������=�uP�N��Ц��I�l�1��O����p3XR<��_ʃ��U?�"��wWt��JGT6Q�93w"���J�)?Վv
��o�zZ҉� %������4�V�P��̳YмI?(�t�i@�������ұ��\/M#��~�b�����P�Ia�o[�|�{�e�K�O��'w�B�c�V��!�[��i��W���J��V��i] ��Ą��R$����$�.��7���bh���X��y��3���c�9��yg��&��ab2�0�q�9[
 	h�K�-gWJ�ʤ��n���B��P��Q��/R�gl'�HU}�<\=��f�ɫ���8zbH朚x�l��/W2:c��M	ͧ�
�lV����| jhK��lӶ�+�J�Լ[ZYQ��B��Zu��R�vc���۽2���������;sw�?��zY�;R��D��Y���
HY�_��ѯ"���Iȱ�}�u��XR@�C5�F(�n���ĽQ!�Q��"��aID��#�O��&R�{˫iB��\y��&t�I@����� �����1�y���6o0+�YU$�����	S���]ra8p�y1�yZ��6�^�s�@��POe�H^SR��� ����d�F���C��x�vN�M��CH���%��0��!�3�A���Z�H�s��l�o����4��ӷ��b��V_�f������⟆OOjܷˎ(��8NFƷ��k�T?�7�G]W��	w*m,�<��w�����4.��.� U����a�Ń�!߿c�1⮹�m﫥㌄�:6~zTv٪�z�����&a1�Q>%�� ˃o������I^�B�8��CB�1ɤ,�)�����O����:�4j���24>dGN��_����̢���0�;f/��$��١_����_�@����J�ۗm�v�5`���E�M�%�:���[۔�9'"��
��V�}4
�.p�0e�O��lUK��~M�uB�3�zαf<X:* @2z'����wߘ
����C�z�/U֔�p�l�����MPt(P�!��e:����b����d�ݼ<������Sr��[̏�%��G �LȎ�5n��bh�瞌⽿��~L"�6��)��׈�z�1o漢�$��� p���(>^���6�lY�z��eHy�ql�,�˫i6��捺��4.(3	��S��;Q�cH��1s�[riG>�����=ҹ���Q���c�N���lС�H��%�M��>60G��:����hW	�!Ê�=嚽RȊoѽ�>/Q���/��,����)�L+�K�ǌ]�57������%۞�[¤�F�IօKs}�J���̲�C�ޏ�!����0�[
���je*\X�GL����� $��u��� �p�}ƽ�����Lp�~�p�=z�cf|��N�H�#K�!U��4s2K:eZ�����G��k���%k�7�g['-�C����ij���'��{| �J�x�g�MM�!���lQ�rkup��6���ɩ%c0��xʪ��Ln���4��^xR�1JVA��A(uV+�׾�w��$�Tpl�O�:ў�p���W�T���_���P��p�]�>A�)�5��=D�����A�U��	�b��POkB�=������a�j1��[��gzp-�~!P
QLo���l��_���R:�E�4Db;nG:?�ۍ}��KE˪
�cl�JֱqK�1��398�K"`b���H-�m�C��Vl]������;h�<�ca�iD���`��DFesT�⏜��> w��`�����U;��`�g��%��\�*��N3�����*�	���i��9d|x:ϦX��}���Z�J��C�ҡ�!�)�_vAM�kR����d��z���zB�SH��N"462��s��(9��U�v�����������\��oL;�.=a�>|������c���� ���U��ôQ�&�8�*{^k�'�jzT�!�OC�U񆊑Vq�UQ�X^��'Uj��ة<���ズu㚴�^U�g�M?�QS`��tû���N�[�sʣ1�3s���(�{���|����b�����O��0�z�U�{���a����ٲ�����B�w��P-��a��@��z�����&���.���V��;�wъ�K<5�WԩQ��?�b�n+I�m��GV"��o��pG�w*!O:������p=e�S�S�C��5����:H���Ն������=q� [�i�m�(Wme)m����HpP�j2��+�J�Q��Ү�0��*}�i�JE��JťEVm�#"[�/ ���P��r�����[�(I��7o�M�����1��ފ�`4J����9!��L�C�{��hm
W���!��ћ�V�� C�5�k�����Ͳ����C��5��bWJ�����0�����L���Ζ,$Rc��_����Y����#s:MK
[�'������]��Åɽ��>�{��u�h�:�φ݉AX��9i�=82��e��$,�8��N�6w�F�ݴ	ZL���l�O���թy~Y4?C�<T�e� b��!9�����r�9o"�~��ѝE���kl'�@��'[-4��R-=�ِ���tN��:��t���c��,�S�k\Ryt])��S �;ze�{��hjbSE]D�� ��6(�]������,�,L���v�|���gF�мR:�������u��b4���|/��4�`⤆� �t��!�����|)�Grx����f>gU���% %��������QM��o�� �9��g�Q	v���Ng�y��u�'�X;�#�^�j������%ca|����ǦQ.b�oLH8�w"���q��h�#�jv�>�������ݓvA^�T��^*°�3��j��A�GJ�������!e��ׄ�����B�F�d.*�S>�W�C@cO�C�׷���5�v'�7�%4]��o�!��d�ܒz�JL�s�<<}��;x�����t��W4HۇL�	�_s�S{�� �4��o��|#Yh����Z�٧�
ؠ��"�<���_�����*���<1fE��˚�!epNs$'�÷_6fk�\��y���X?Q��CC��~����ġxS�1{�m�5��[5��?,.9)������嬽u���q�����|��7�C@({�4[U���(r(�ޡ>�[X��gQ�+rZ&o�]�NNƖGR��0�>�ɉ����	;��w��/��?̡��k� �Wz>����T6æ�7�q����P���ʗ����^�ȁ_�z���
�:�A6Ɍ"����S���4pC�Q#��$y��������Vs�<�I9VW��_�����	�%Ph����x��*��gu{���w�!>��G�)_��OQ޸AH�*�Uf`�Y�p�Z�08a�Y��x�z�&������v����@�Uq�<�š���0��%�o�$���!�ٮ��#Y�����B�#��(�F���K&�9�0jn�.�4I�$,(�e=:��^[a�ù����"R^�K6k�+f�<�lf�V��N�!�1�K*����"�P9W�u�'G~�Cjݼk��Cŧ���j�#z��1�}�����x@]@"�ut(��u,Pp�*��br�~.�&��F6��i% �.��P�i��\'��R*��������/��H~W+�E�H=7�@�fĀL�7��ӛ����s��rXm�hN��˹�z9mak���������E��7��`��õ���E�ysQsU��k�|J�-=.&�A��.~<gQ�� lH�Ƥ^8L̀���͆�9����"h˱�.�ʉ�ھ����Bc1!�o����k���3H^��2S��S%���U��������;n
��S6:���f��A�~���M#t9��hiM�:i+U��/�/|�D�<f���ܱ�ȑ��>4��!?}�:�tf*ѳ"P��|?��]���"Ͻ+Yh������1���e���K�k�O�L�(5^��v��8:t/�}�O/o}��a��~~g�<���.=C�x��YlI6�!�����3@~���:�a2��vB���9�_�_\̙H`�(EC(yJ�0Hv�(������l;AiB���MQ���]�<���0�V÷{v����� 	ͯI�O-�B��Iġx󜭩crJ�+I��ǐ�I�I��(֐L	�Ϭ��
��KP/�Y[��Տ�H�<��1r�B!�^`�4B���8��ul'e��0�v��RMFN���eg$��魙��̮�����7Q���b�S�k�����q�m��{���]���Y�2°��a�|IŸ�*�����`����:wQ*i��}�%�Z�|Ɖ�3�����.=��_��Mp�P�������q����V͎ˠ�
��2���Z,<��] ����tko�[�]����9����:���o�ڞ�1��]`�V�W�Ċ�'�N�n���Ԅ_��Z��y	���S����ob.ob��A"���qB����v��K&�k
?�)͡XB
��n����}+s%�Y�y�:��G�����d5��ի����-RY�)0���;�F�r �Yu'�p��l*����?�����s��R���f��ǎ*��T�qTs
���}og�S��~�T�X+�|>��/i&�Sb>�A������(��N5��m��/�7]n��>�����,�RR��dA͔�w+�díHH�ܫ{������K�ԣ$V�r��)򡃩Wv�����!��V83�l�8-7�K6�Zg'��Q�K�a(���?�dz���T�E籶��Δ}�(gan��_+,����+��V�|���.bA���/��[�iŬ�w��t�o��2�׬�H�^Au��0.�pt���Q��!dZ�	D
��P�<�������1���#V���SN��~�p*xj�1��l�>50��H�Vb^�J}�DĂڜ����	&�����H]�V��u����m��f��{��:�������c�%�m�z�є�^|zcU����k��c[2S��ԑ����E�;@Ib/ �GU�n����~�tɶ�|*f�m��5���]�l�q$�.qy	�Ez6�X�aV����B�/�>��7�x��m���)�!�+zy�F52E/�E������*�Յl*�[�(��P���+�A��3��|XN�j}(U0�$�rV�pQ�י��L�%��wϏ5�b�l7Kܓ}²� Փ��ݐ0D��ՙ�9�C�������'i[�f�$?V=B(��P�qJ�H�bI?FZG^��P�U �~����[-|������
����{��X���\�W�}��+\�,�����3Н�K��0*���Ƕ������G{jp��m^�Jn�pt�LI�eY��n��8����M'"f�� h�hĸv�����:,@���"�`sp�Ƒ��Qm�	27.�+[��Ȁ�g��wG�5Is�D��H7�&N��J#��q|���\bJ������!TE�ڿ�7l�*>�TQB[�z�%���w���~��a��cیW��%Ȝ�Ϗ�l=M3(R�y* �J��6M����G�����F��Z!�D�,����]�=�N��]�+,�Z��i܅�fZ����)�nǸ�Y����YJ�9}Ң�B�Ԥ�8<&�i$_ 8P�6Zq�����t�gzK�kN{�͸�A���c^w����Qd4i��d$��Xo�9硍��d֣v����!��"_b,U*s�V���d�3r�<����T�xbMy�i`(GJq|�w�r�s#Z��c����1�޼�Vl
�G�*��>�����8U� \�TA��dݽ�����-�|r+?IC���why��R:*�bH[��.���Lth"%����´�C�u�ڒH�f�����?�)��ߥc�'�����{����
}�����Fq�SFne�OP#u��j�s�~�]�5Vǧ��'~�Vy �0q��L��ghM��Mm���B��0��zP�{�z�$%�w����K=ס����N.E��s$�ڷ8�!�d����!P(68������n������+,�EFkyXά9�����StaVr��>$��u����C���ؘt���ۉ\�m?!�
� ���籃U"��;���ӳ�0�����t34�d8L�u�:G�(�H�{�B<�����I��o$�~�䌹�I�EF�y8F՝5�O��{#��7��X�Y����_t��g)�?J��
HC_�p�����j4^�^�а0��wH+����U���	]���O��;8��C�ӷ0�>��v�ϯv�s���xA�hU�=����=+��$�\�}Mh��c����
�}8�����w}�T���u�"���b`b��̩����Dl��@.!L��T�P0Q�3}�;)�zDB�Jx�}CkpR�\_I�T@�~xH��M:�h�T����(��\�ڕ�ì���֟5�1J&M`l׎�_/���7Q|!5]�ŧ�)����򰇴�OuY�Bֱ�?�I�Tx�I�����B.�g��c�� M[����i�be�$�jGrU�Z�>�<���u/�ZCk�]���ggZ��>����g��}���LJ�#uj��]��(��ݸ����@q�97�H��к��̴�T�Gӆ\�Ɍ��]�=�r�w0k�U�M|ԑ"d�SϠ���y>����<�4��[
��M0@������>�9,�=�������JP����d�<�y��@2����Ч��ێR��X��'ԣC�m��RV�%� 
��KN�U�)����M�*+/[0���/�O����3e�Z���MX�W�r`�v3�)h�C�FWVj�
��d�M��G{/�CVc���"�OW��9�rk�zm�8<�������R�(���]&�+!s��J�N��؅9��EXhrU�]m���Q�ѣ怳 z�M"��>y��j`M����y����N:G���F1��""���/>MO�$���0����O۝�PAO:�!F��+�1ǎ��U��S��a=����;�B��^rO�������L��	�-�h����=�o��/0�?}J��t��`
���!]�*�q��{�Ū�,U��ʟ}E'�IvX���x��q��U�y��%����-t�b�sES����5NTE`� +/BW"&��a�����,����l�=V9�O���]<�RqJ�S�������ED��	I������i����*�pÄC�Q�Ґ� ˪ؙ��O�S8����hq��������8�2������<+M��P���N])H���^��Pm�������0�Ĭ��Ҏ�e�� �c��>p弻Mz������n`k�z̽��fjճ@I����e�Q}�ۻ�������P#�LK��z3��\�q���8���4��F��D�N�׬�L��x/�4c�{�ߊV�aШ���G!��9��[A4��)�[9�i[q�m�(����1��`f,���(k)ټY���ʀ�}s����3�ҹDtvW	R9	-ӓj*a�7Z��
u��z_7S!����.�� I��뎸me����-L�kp7m�`|�.nO|���!	��F�`OzҼ�7�WM�K�;&�#:��o����p�r�wܜ���55�BS�Q�w)�.6�ϝ��F��f����Fʾ �ޑ�I�m��B��h��;=�61�pԵ�;�@�џ.�37�ۚ��z�Uׄ ���zp��p�eyR�3ĝ���5��-��Q�.S�<T��׏<<��	��`Ar/B��XSF��*�C�ҳ�裒۝��H�����I̩��>i9%�Ї��Ɛ��`F����2��ͻ,�}�R)�;<��=���nK�j�r�r�v���Z�v-Ѡilp�I~�t�'�q͠����w�sQ]&+%����3�=�ۮ��U���{C�oS��6B��~H�\
�NSj�:�H[����q[R����!;��Y�K���,Q�v�;�6��q �*hK�Ĭ�����0Iy�@%��HB�&��z�:B-�&yc�xdf�z	��&4�i�zYE|����Z�[���ՠ5:C�k�75���x#C�����֘�V��?�p�J�ۍ�R�&����w3���=��F-���6ֿ)�z���jJ�������֤�\�F�u ��`E�%�gob�(���y���xk��E���ی�P�QP�/��Mn��ɗXZ���Y��n�w��~Ꜻ6?�U��_�=�$έ���nΔ��$l���Lb�G�+|��{�+Gs�
uÄ����'��-�Dvb�^c�ZA;W�i���Zwְ*[hJ��u��5 �ٙ{��ǯ���n���2	�<V�^	N����~�,��ed@�Q�><�߆��p|�b6�9<�w��#=B�?�����C7N2�^8�I��M�|��}����\>�^Ă�}jŝ<�C������ԁbߪ�I��(\�Zcn�
�H���㋏B'�ڕ�#�Q�Q�e��_���3>���-�5�V%���,xY��sk��)!��כj�>�Pz%��4N��B���'!�0���*\n�m��Z��P���l(8x���-f�
�((�8�Z���*���
Ȃ|>�(��ߦ�X)Ô���?��ߋ���2;����^��_W�YdG�Q�]v,�N4ke��4O�Z9,^�C������I"��do�������~[��AX4d&��ka,ȳ�,�m%eJ���f���+�j�_�E��%��'�@�-�Ac^�l���B�����ʹ�%]���!�7�CXg�]5����z�=Wt<���~�R�u��wȹ�C(���7�"2�w�Ui��M@�Ȕ��V��<����V%��i�/e��;��܃�j��{i����Z����Zҵ�#˕]v�Q㱚xo���9�A�t�@ŜQ��B�Pj����
@KҪV�ɅE���b_5�t��mT������]��J�}���V�v�B"*���y�H���	x�r�r�<�����Mj���`��VI��(������/#��)k���r�,,�p����D/�?@�!8�����	�����1u�k㊘�$H�gC�ZeyG�rH1-��Ӕ�GϞǵ�^3� `֦Uv\�]�`>��ʽ�t̦�&��2�/�d��4	�R�o�΍�/�Q�݃k��\�N&��2��H�H-�~l)�Rܧ�|Y�
�=�,�.Jm���TaZ�����F S�@�精0!���"��&P�����8�^����h*)o�ؘ{&�3v?j��5waJR�j�p�ǉ��.�4Y�d�� �a-Ϥ���2p��`�:��=�۹ǒ�qZ4z�r=��Gt0`���)�����-��>p��{}V����9��51���SlF�ٲ
��̋a��A(d3oSPv��ә��r4w"���1�~Z��%��Z�ӷ�h�,�ζL'�y�~'�{��@�+�1�dM�+$1�5��vP���G�S��Rߨ��*�$�p����lz��Z���#K#U��\���� ��I�a9T�"D�m�%�m��\Juw
���;9!7B��V��Yc�l�I��p�
�i��9����g��*���B��d�0���kUm��_�������I	Ϧ���ޤw�2M&�!$�U ;T�A�@>n�;V�A.���gݤ�==x�f��IL�NK��i��.@;.�=y�:���CR�����������!4��`a�M憛�Y*ϗ��X���UM���6N�t���NI�������V��q\,��3̲��ʼ�;=W*��2��|z����v��F0�g�SGL���E��	b7x�/VV�fY'q=�}��D+��`SԱH�Pvº6�545�y��WX����
z�˯�x8'�st4�I6�?A��  ��lT�DI6��zM7&�^-��ʺ��3���Rg��N����T��E����O��{�����c��2N���w�H*d�f[ltR�}A#M�jb�S�0���[qu*Zc�܈F�p�2��ٚ�/�X�x�E�[���_�xt .P�A�T[x���P @)��}�TSK�}���Wg�U�<$S%���+��XOe"p�C2��8���ּ�� �Ƭӭ�Pce��zM��~�0��RӮdX��xĘܮ�s'��U�k��Z��ɨ�9�C� �w�S�>��u�+y���t�w������;%�# .F%�s����cߞ{���v!4���d���|>�) X2��#K"�d.a�fh�t���2m4M�Ŭݎ����^�����	�3Τ�i��b�����.tω56I_�ꍢcؖ+�����A�ڗ�P6�����֓���
l%ݔ�b�!��T�0��e>�A�JU�\a�|d�ǋ\o�|;!�
�]�:����6c|�nVGƢ�!�ӨTA��E�y�����:���Scc�⼺E}k���"Ý��ƫy�m�8EK R��R�+�]ȨT�ۀ����K�����'}Vl,�m�+���e����m�N�$��Z9�����H�<�=��2��q�ZP����z�"jW�ev��5({b)��l�%7��3y�cYq�g�ҭ�J���:�é��b�{5̤��df[� �k�*&���^�[���}�=��iQ���,�í�"#��rS����!e�\[�'��E�"֦c��']��X$�o��4��v���9�!=�Zhl��|vm���<�|f�=<�ϵ�L���	���1m6��N�V�zn%��r�KYX�ʥu*�n�1�O;K��tl0���U��ׅ]�*��Ѩ���E�o�xa��IA�tE��	'�����k�Dh��|���w@�k3.3�p���Ǒ��a��M�fp,,��?7�n)�4Лԭ5>ːP�s ��vDl烞avq�v�o����`�j�R�q��P���ӊ0rq���� L9��>8��/i=�: s�?��9�SL�W~�K��y}S�}Ğ�$ѻn��;�
+R"��[T��]�R���hY_/���k�o}��fIC�����$X����`���j�T&���<�	`�Z�vxĆ#�NPO-1�1Yu�%���*ߧ�}����̺ϊ �y���P�L'gsi[tA0�GKn�9/�6��o�ptri�)f��T��I~<cywF��>@���|R�q]{�?f/ \�_5���g��B$�K�#{��Y�W�L�k�4ޣ��wg���i���깺4�%�0T�je��ը��ֈ����ƧW
�y�2� ��Q��Y��ҝ�j��rI��=n���UB(�#���V
=_������:\�(M���l�5��Wo&��T����ڮwOb'6��*�c�iY�����jG)�aH��n�!j���r��0�U+�Ov������b�U1mϞ
�ZXf�=:#1�'�t
{�@�R�������_,߁nX��M۬�MhL'E��lnM��WK0;%ff6=W!�1�F�c"e0Vз��Ffҥ���g1�g;�M����M�Q�����h]��Z�8�S����r�����<�ag����za��J��@��#SZ�W�;� ��_@��_Խ���6������bsOhWq��sw��.(n.�S�wЎ��!�ObBgy�3{H3E�H�Xc��9N��+NHr+zE���1��RȚc�𧜑uzU~�ٯ�t��' CO-�q�ڶh������V3a�3h'U�]�I��P�/���!z<C(��+�is�Թ\B�S��L����/�(������5LD�M$�ͽx$h���	^�SSP���A�qk�}�5��قb_�u�7��11P4��8���پ�A�Uk�,IX��H�����s�E��ib�t���2��Ǆ�d�R�����tiH�^�@�ˬ�H��Ld��$�
�6o�j�����O�<�%�:�܍y�[s���m �>:��:m��|Xر�.XC�+yA��x���e��4='f��T�~��m�!�t֠f�>{��~�Z���q�l�U���yj���z�x~e��|R��L����Q�>Q�.�#vK/���~�n[ewE�nwq\��2�%B��+� �&�nvM��yB����yW'udR�Fu y���t�DthnuUO�OĮ�b֛@�2q��j��o�32dL�7֞>�����O�7�?_�&�<��+#_$i�C��/�{�@j��uyEO�^P�=v�H��)� Xc���4{��{��>���F��>1d�l�jN��b��M`�[o�.�l���"��4=5������A��ܠ̙��琕���]��c�2��	Fd`o����F-gx�Tm����L�M�+��ڿre!�8D��p��cQ4��� �(/4�'��$�� �v�f�d~�<�o4�C��|�
4�e�������|�c3.@���shpy"2l�����G��+�ܤ��`I��χv��� �O-3sbfSdڎ��Wr��D".'C1W柄35�=�g٨��e��Y�G�_C\�rU;�|>���# q��bKee3����u�#?���<���6���~�)��M�co%F�@�v��;A/�ct�Y��ꩀ?�X���@�������u���XX�膈��&A�d�p&�l��ț 
�t
fL�1�i��o*�E�S���� �Lj�Ś=Dkܥ���<����M��m���΃��n?=L�a�I��NI����GY"�ϻ��
�Z���y��)������,�8B.{P�a:P�@�뽩M�Sw��aQ��ms��[��tc��z�,���V:�h�Kz�#:��=d�$G�y���>��X��,���?-m������$:��r�,�Wj���TI_���`��n�$��T�6�����>4D(�S�=TL��M�uX�>����Uf�ϼ���� M�R�1�@�ӑ�;�Hl����Au�����t=ʮULڶoų�a��Wg�3��~B�R�T�`}�떞�^'���8q'���G\��k(��l�L#��8,sg�!��!iqw��1���mT3����t�İf���C�H�%�!�'%;�������]�ѻ?�u����UӴ;ЇmSY��h�%�#�_c�6�%��.y�L��!E�F��l���:T1ѱ�?�,��73Z�tFW�6�^����=�w^{���ٞ�D*y���C�`��K�Mc�_�Y
v�ε��_`O#7ןZ@$X}����vp����
�ۣ�U��ݴ���7_ߧzԐ���&	82��$?v���f3�^�(��_G(��z�cs��#�栈����/�Y_Mܨ��]wl`�)�0�xe���dF\����]OF.%��=� ��ܠ��ߞ{�ѓ�����Q5�F��V��F�v��n�YQz 'i;C��`+D��0$���#�j�
}U�'��Q��% �wd�M��oBdP��J+){3�P���&����`U�����wG���ۗ_���W���Zr?�AX�$�e�>p�j$�J�į��%���loa�.���t�� �x� �� ��J�Ma��Q'3:r�3�r
�y#��-�b�]�Hu^�7t��]c�	q8��]���(�s�7ɕaC�������Z$"��n~�o{NCJkH���Q�� �e�o�U�L��&�Q��[��o>z$���[��4jU#ؚUa{�ȏI,���'��#��?x��z�`T���)=j��Sv���=�vs����0�8[Z�%�>��s)Dvbݧ��B�xgL�1p@ǌ-���\�Ȋ������%X<K`��"�� �𘃟x��lxy�OH���� ���z-�4pny��(�a|��ƇZna_%�]FSv�~CP%z��2ũgA��D�4w�K�LϜ�D9��|�P�]:�9��}A@I+"-��%4�-y��:V�QI�۬�B:��=+�H�`�xQx��M�naӅ`kWp����EX�5$�5�I� �\�D������m%��r�����]�P&��w�L����MrO C��SӬZ�r���-!p��	}>^b]"�?~wL��4���x�%����zS��ʞ�rk�0�Qw�&��d�7����9��F�
n1�
I.��b�K�����:?��V�x~���{��"�|YJ��	�k��iB/�����h�������ێ�E*���?
���△�$s2�%������88�W�D�^��83��2_Z�
ރх�Ň�ŷU�pʼ�]vjb,�Dn�k�|Hi7"�K��<0k��II��TG�H����:M�݂�v�k�&��s�J!\��HS(O��``˝��*��������A�e��$=.���`OYvW-������;�ߌE�����j�V��ࠣ0�A��D|�N�ޒ���m(�+�����>G��,�c��e-��9vN�]b�:j\�f��є�q�w]�x�\�rn"�8CR{�E��V�4*��{ȅ��� i�]��qJ��F���t!e��b���m�O�Ưo���%���I}�09~-�������8�.y8gW�ЍR�.�__;��]sRVw�����}��z�Xo���q�+}�')�O^,VT�$�@���<ׯ�_*R������?��_:�p7:-K��<V�a�p싫���E3d):Hf���ܝM�����@�~GC!RQ���A_4���(�ygЉ�\sP(5#��.����<��c��!�]���������ƭw����z���
���ڶ}9Y'u�@�FOA��<�+�)�.2��$�:#a7|�>����\��H|�T�w��!����@��"=[k�v2t��|�^Vs�Z�Fm���7"0<�2��Հ��.e��A�DQ�6���Jȩq���������|��/�W��\��5W~u�����<H�iF����n#���Q'� �L��� Bkw�Yw�!����Ce�j _�g�����K���F�z�Y���0�1� 	�>�׭IBl�FiPm��Z5�fE5u�5�+-R�e�E2�1!/�r6Qǰ-_V�m&~�F��$���ƣ�-4˗��ӌ����G���v���?����
���F������}Y<|Qo�>/ݣ*t�����u��M#�hJ�b �z_�O�R�n�xo�geP�������*?u�Ki&G�ˣ�$�G���r{&��oѕ������_w���9������_�)E����@ʾVԩ+fJ�=?}�	�;; {-Kaw�{0�m	*B7�4~z�=��ZN��ʅ`��_r��]O�R���?F&���\:8}�s��Qr�Rj�A�2��sr:VZ[�38����8yG(_[8�.�	��m�������!����*�ts�ʆ̊��:�1hu�u�qK�>����'�g�?t�����cR��<pە�~V6�iwe�s�˚ᭊ�.3��`I
�*{�d�Tu�Q� �2���<�Ow%�>d�<�א�f!�#n�bK�&D�!�==l� `�7�^#�m`��(������_���TWM��Y!~�y^=�p~.<h����w���sX��ݬ䗟=�3���������T�}᭓؈b!?6UL��ށ�Y�鴊�h���!�рLIS&���H%}!�\n	�Rߌ�e	����솃�Ǟ�p4q^UR@6���z�
&�l��
��y1UB���?�pẂ���fjЯFx�˻��mç�6קP��_9���f(`<���؀�rc��
���d
;�aUqjckM��
�K���ޏ!ګ���pl4F夏%�Uځ*��#����_l�r{�hO���W�𕮢�����u���<��O;U� c;as_ߐ�<�:��n?̦�_�z{�zX�� �)o�\\a�9�3���lY���_�C.?�ڜ]D--��\k���S4m�֖��Q���r8L�\�jA�c�
�A,flH�O�N�)�$�c�y].��{��0WV�̇�G��Q�6(6k�2 #��.��v�(W�A>Z����J�A�/�%�;�1¾��Q�Z
L��]��!*rI�^=Ԥ�	�w����f��-���p�����B�?��'=�1l�O6�@����|cW�.�Fڣ�U�H~��ДЅ �����������\C?��M��Nf_�/������d�U��T���U�F�)4p�>�B��o蝭P9�����I޷/��}ϰ�(��=���	ь���8�Y@���I��g
��$�Z�=f[xxDڎr�+��쮗�/h�H��Nu��-\�?������%W��k$�t�*l��x�F'��{o�w�3 �ڶ���Z�6�_��`�����7G0���m5Ҟ���46��	��i�J��!���<یq�s)ʦ&�ݩ�J�J���Ȋ�LYp����o<U ����R�S��3(+���d��H�;�v@�<�����Ċ)��o��%xL����0������ �K����h��z0v�Ϥ�FՉ��)�%H�߄׾���~��Hz�c��g������g�,����5>����*e$*�tUG����w�i���]㉑�����f��UȲ�Z�$nQ�YQ��ȣ?�
gH8��m~�4`�f��?�k��v�rp��ѣ��2K��z�$��1�h锩��T���uL��d��f��rU���[�D��fH���lQ.�I�)DVե�+0ѽM�^K�����:�!Lgp���t8Za�y0�}�m�kD�B��U6qq���M��d��T�>P��ˌ��]�FA�;�5�31+?�������/����tS��&T������u�Ǆ)<�GP˽�B_������m�OJ�;'�6� ��	��#O	Z�3�:���X((v�)O�O��$q5�>řR����V�8ӚGDEjG:;%��,��i*(ʝT��ꢛ>�H��>(���<�_� �|�L�/�,�.�m٬Kwo_ʵ�^����<�g���v�{ϴʦ����g��ϪI�I{V�!�?)z,@����(��Ț�o	g�ЗL_)y�r��a��� H��m���Q�IS *�-��AIO���}�3��4��Q0u:9d�s��@Y�JoY���	q��/�B���Z�������F����1X��;��w'a}��	�����[e�-�}1؃Eo��~���=���R{Fq#s��V�90oe�;Q�Pb��3�Kw�6��[�SboBL,�tx�O&���8�n&3��>�J�z�#�q3UgXt��iP���[� :3�g� 2����y�5Or����Ȗ��\��KV���c����r%�����B�_�M�^���G=aCHsk�vӘ��C������02o�um#�!��������Q�ƓzH�g���N�mɻb�8��3� ���ms CLmR�F��f�\Kj�o�Y)�3d�ƫ�m5A����&����$�/��(��]�!)��zkw�l*6����r�7^�a5%��kON���lH0ZS�D�lt(��Z8u]�i�u#)`��Q�W5�7	H\yzY��_��I��l��1;K�&�%b�̡a���}5rU9o����A�H���8�����bU�r�3��Ey��9u~Q��0�l��f��_R�V�O���l�3CQ����v�G�.8Mm��P��Z�(�d���f^L�&G�V��Ǽ�$�b^p�Vs�kFp��yOII�4�[w�sE�F�-X�����o v�����B��Oޥ�3�,�����x-EI`�7�!�o�H��� 8/�5�L�%�$�A}%>���4�,�n�%kZ�����dz�|-�Ub0��E�]A�aDa�h�;~�#��G�bL#����t5�U���Iqgh���u���4.r�w%��(�ƒ+���%�/����R[,S���"�T0���2jVB;�L���ophu�)^�}�R�=�R���l��F�@L��*��
�0�_�+8�����W�Ί������m06�ޫu��ui#p�e���4��j�.ʩ�����X:��+�q�X H������I롁U� X�ۈ�.l2pL_6����ُ�3i�2)�.�83�`���U�۱J J�á|��e���Ѭ�yR�$R�՘��C�����`�KtD�a+].����:�/Ofb��n7������6���OUg?S��E�g�m_�K�����;�����e~����~��Ķ�L4�)}erzG=LB�_<�x�O^��I�HB�Z��im\ۏ��!��W ��,�Y �@�#f��;ٮ�@�09#�j_�\F��}��a�(	ލ ,M�y�(�]���u"_,�]�U�1j�h��;�k=�W>�u�E$����}��AA�=	 ��𦛚r,�:2��W^;���(c�
�@m��<<nM��M{l�*�V=t����+�r��&��A)nԫ��ͧ'����2t�G��)wn.$]�,��Ī1���T<����iǨ7����!���^\Ե�G�����7H�~.�``�����u����n�i�)f�
y�I��|���
E�uL���Yưe�&�j��v��\1^x��ܟ��E@������wz�J�#��+��ѮAlpb�O:#<�S9W�FLA����L��k/�7�n�%�VccD�?|�`�Q�1��z_;���#3������t~�:Bk�j��s���Mn�o��8㼤�����v;s�6_^K��"�4�}�!	�Q9��ؼ���u�����v���z�o��3�mV��P؛%����8�+$+����[aK�����Oe��v^�gH�3Y��K�L/D��l�U^���c��k���%�YGĔ��/juF��o�,,��1�o��^;�~#/������˟�_�1�&t˵��)m4(n&р�mKUy�?NU��c�.be��m$��r*�[��3���PB����v�M�%�c�	��2S��7��� /�{�+/��V������	6��$"}�P��G=�3��䳂^K��U�
	qO↠�༷�����CS	��Qf��+�N�m� �6.g�mGs�;�5~�J��]�Zgܭ����t"��ƻ�CS,�'�;�51	��Ϧ�$��'ИM2�FK�8�W���fi�&���~5�}��_r�	���LrE�n�#��X.9��ځ��0�δ�����h�6y�,�ʔR��t@vP�]�E�-~�&^�0�E, |�ŻS#�F��hn��{�C��������i�5h�ʈ�Fv�{�[�q�<�3��o��@i%�z�=E:R�0��c�	��3���
��jڎ�^$8����i�YN�B�"f�x��u�������a�ᔺ��i�����hP� �hDE�*qρe���8\<wz�m\> $5��ѷ�x|/������pq��T�I�,x�/��(. DP9ߚ[z�u�R0`�L�������`hP�Λ�0	�KtV�zQ�~~�&��2y�룎�`Rvq�6/�� y�Z����|º��` @n�����~!������;|;b+�f1��p��u-�N�)��v�Aw�P�i���.p����1I��X�=�s�w��L$�u��As'�|�>W����~	�� E��ӲxqeRW��_�-t�D�L�B"�xD#!��]��r��O�G5S�9&���2����vF�o*A�ڭe�f��5���T���h?��t�ޢz�F&&*��4|*@-8N�Wv�,؁�MG�8�ȗ��5���>Q�8>��f��,"� ��V�����դG���y����������N�)���r�u"�'�ʐT,�%ұϑ�{�ʺ�~�Y�Kv�+�<	�h����<�����'�E��أ�Cg< &������E��a4߃U�A�J#_Zg��d~:y�3Mv�*������?��=�ಗ~���a���[�S���YdC�u������/�F��M���h_��Z�W�c�	K��2kY.DsƧ.����b��7b:��c�|S���g��*(S�#9�����{(�\E��lv��L��'��- �]�Š��ihs3g/~a�D[�+�҅�T��<u��1LT����
�9�������\<� _�����]����
U�~z!r�����q�<�j(A�������,�0��!��;�?�\�	�@<-u谬&��I�\K����[�rL#�bW'�VNiޞ3���V::z;fkRU���C��eڋ�C�W<w�)"ݞN:�����������B5��T;Y�� �H��P��^HnIe���|�?d/'2�^����
|�8��8�h����h�1-�rm�uMD�k�*�0c,di ��:U��q�L�QP3�;�AiɄُ��5�����B�L�م�
SfdO�g��fF1WH!�Mv7s�L�����ɫ�x�'Re�dQ�@-n�����MdE��)��Dp1��=%"2��\j��o<ny�U�p��#�ԐG&j�	\"��]�C�[�1�!��U���گ�̈́X*qJ}8v�]��.��-g�:��8X(�E��k��*	�xh1�Q���oie�s���{��9�<&�������)x�b���w�8F+�Y�$*SȠ-_fkn9��炍|��t|'���C�t!F�ݐ�ϲ�`��C��u��4���%�o��2,{(ӳ�qR�ā�|�S��M++����XA��"�Hљ8Y�O�E�͗;��tT�Xp�	�s�3����`{h;���$�QK��H%�=��wF*��P*�u���

���Eљ�IP%���W){6�u��e>����r���ыvw�Վ6���л���	c'D��B�n��>�=++)Ա^r��Ga	�	��e��$!M�t p����:��vW�X���w�ڦ�\��@�59�� �}���B5�[�jh|U >5��Z
���8��߅�"G�՘}36vy.I�x;B��	r���d�;)`G��L�c<�a
#d��������W�皪��ܗ�V�����H��� ô��±��'�Z��R���\�Z�����?,��
s7���8ؙ�%f�����POXd~x�'���XB�%��4bm"����&{X$�>ζ*xa�~VF�t8���o��rm{�Y�U|%#�����r�}=�X-���paO���5i!\�[ce%��Q�a�\ߖS����e)�9��I�=��"�iOq�ʑP�m�1�!N�S�$3P=Z���I�hT��Iu�a������`0r'����D��$�l��0�˻�\�ȿ�3V|���\7������������V%�;�'#N�W�"����^�U�5���W�O����>V�q�;�3��}a[�_���Px�唀�E�T��
�1ZZ̴Wv!� �H����x����,�'�'?�.��9H��P�z����
���>+��Ƿ_@����sf��� 8�eT�����2����@^��G�s�;O����s����G�fF����\�\�qR?���nqȡ��雭;m�o�b����������N��F�3`Wu�R�PX~Ǔ�WS٦���ى ��:�&�;���=�]i���z�VtY��|P +6m��T��Gq��&�\mN��X��Y|y��*��pe��o">g��!�Kn�g�y�����tݫ����|L�{B��T���o�z����D��L��!#��8e�a����΂%�ɱ51G��h����Li�ǝ$	=q�6'���-�h`m-�3|�Fd\xkN;I�F��:�
t'<!nvs��:����\a��<�kU	�<R�cG� �Gz����M3A�f����ں��8�J�%:�������n�w>X�hɾO��/`c`�E��wH���ܦ�{3�GS^���r#�2�-I�Q�_
mq�LE�n"��Np����mWl�1�'��h��^�4X ��eݐ��WN3݆rx��;	J3�2�ek��H!^�ķ�ASˣ��G<����c�A�8��ɕ����V�H�A�+]F��zy)�\�K͍�����a�Y %�#�i��v�x���G�+ ���Y�0r�2,��n���v�!y���t�3�'�;�:xka�4�L!�b���Ӻ��;�s�r�$�9G%I�t��_��m��Z<C.=|,��c|C��.���bL�f;`��t�����C��=�����
(�
�	����m��fpd�J=�	�.ؖw����w���*�MΘVM�2%���XP�5��友��v���4����8>J~l�/]8>��W �4�!$��p�:��ѡy\m� :�:1�vvq�Y�L�U�~��O�|�{�J^�_�Ш��6+���p֛
w�U�X6���랼M���'h�������L�LF1���z����(#g�֮��B��]��J>���R�v�3��T�8bk�g)	��x�hQ��6z��
7�K����C����0�!���y�֕j�'�++�f�bS�ѽˈ�>��]IB�P
{�{�˝s�i�)Ų�	Sǧ�����)D훽�Cl
�gpɸ�6AП[-�ӂl	�7��q�S9x�E���!�i18}Yi��!���zRY����-�>�U��;f��Ө����{��ɼ])s/՜�S"��{	���R�//���,mOʱ}���~Յ�``����س�l,6@��7@=�V�����:�J��~��2@�������Vo�C�|}�?h� `�䦫�Mw>��d��k��<F�]�B`��OR�v�6)�%����>�i����9JhNA��lĜ>Ӵ�P4/s�ع�G��GW��NZ�ô���DȊ|�j���������D�Z@�H�(Y��nqHe�yi���$J��R���2�N��?���y���Ɣ��`�M����l�;�Ѵ��浟�0�;���"C�?aݮ`�I��|�Vʋ�>N&�ݶC]'�����0�a`�oCW֬���u�Z�y����ˆ]�@4�`�7v���8x����絍Kͅ�B�:p_Å\�#��4�m���t���T.k(a<��=��9x{��"������v�2m���H=^k�7/�6CɄ����L�o>������ "$YJ�u	[����I�J�3�O��"|�,e8{�t�<��}'��oZk�H?j�i�q��߃����|���0�-�ϒ��S����;���)枞(-W��b�X9�������&}���d�b$�-��S���;亶�]a�U22)����5��>�C"��7#�W��+����k�y4̦Q��M�
:�T��.m#���)����\+:{=B�l��oz�¦��*߅�h����f�?��\6�.Eɼ�cV؅�mȈy�(̥���/��t���~B��F(+VӖ��+Ӑ|k���K&�lş�}�b�}c��fѪD �����%�q��"e+%Y
Qo]d1�*�����E�/ȑP]�4�7������nP��z�i��2�0L���j��mR8gs�4v�p�&X	:,E̝�z8����u�gE�$�*N`�|�FFS�:�����@��{�f�di�v��,��R���t�ͼ���DC�_O�E�C��x��B��D�(�A��2
����u��5l�r�����/E5��`������õ$�_ %,#�_%��¹���1����#Fah�?�>��+E<� ��p�̯v��!�p�OǸ���,������3����W�7-�nO!�a�R�^?� q���� ���3B�J�ߟ����R��y˥K� p��j�:��
��(�RSQu�Ko}���S3�?����%$�s�OE��l�C�8�P	MX����e%32ƕ��`z!���B�_���F��:@�9|��Dj��	r�0C��ڂ:K��7�dc�T�x�r�k�( .o �).$�CH����9OTjv�˸�V����2&���^Jf�m@�߆4�?������;5�f.�o��/��֝Y� �t��=="I���t��:�y���>{o����|a�VF��+v�f�eD#2���n��vL&��Z�ɃP���&��_�ХX0�
�\�RB��}wK�fMI�jl��c�b
b#��abLA�ChX�뭲��=��~]4�x��Gj��3K�f��PE�]M�dSW)`	0����hOB���L�I�z��k�������g�qL��5[:���� �C
x�h��~,#�x����m�Rc��q��7����Y�~/�����Y��Wy�����J�YPj$����ghǎsR�}�K�o�����_�l������~�TK����X=����q�L7*�l@���9��3�����&^`��]nL1�h^��U�ou�qS����	]�Z�/X��ǺN�.�|Mx�2�+3,T�'�\"��ȏ��#�e}H}g?=�P�ϫ�ʤ�G�`�9��y �7 +�`O5�&����j�����L��^���-������-�c=t%|^PGS2x>�X��ѭ�[��!������J����<���<��[��fW���N�k�)��f��Sd���%s�Y=EJ#D�����
� O�|��:�r0���N�H��X
M�K�R)�n�-�:��$��$��㊢��0s3�]%������6���hj(G��Ņ9mg,@��L�1�c媨y�f奝�~g��W$�(EV�J�7Fc���;�&V�T�RV����Ѫ�p6]��7��A^�B�>R�U "��۴),�t�V�~���CAM��b���E2�����	�d����{V�������.%��F<�����6�O�j�e�]8��g6z�/�Sk}���c:}��v�\U��h���Ķ�}KĒ�p1�2a. � �}��a����Q-�nA��z�Et�,z3� d�sҁ0��C��������L���(zFt�(7n�r.p��Ο���}���ԏ��u����8���!<�Bd�_�x0���=Ѩ���ސ�Чy�E�|�Q�F�Vu0����>��3�P�:��U@�㎧�N,yA��GP����`2|�}���"�2�8�H���Է�Hڴ�zK���h�RD[�g����ݒ�׬��z��M~�/��'��'ɐh�_U�FM�~��$&��� �[mЕ���IM�E���6�oKz^%�ٽI��U���@��7dF����eC��>�{H+�`?>弉e���'\���J�O !�F(�Ԩ6^�g^�����󣒶8t)��*�GhL��	%�ďQ�p�0���K,�u8+��E���WMᣠ`{�J-�UF�Y�5�7�'Қ|�^�����	<�>��f��JB9�)�j��`��#�}�!!��D�\��Du��!%����OU��xU0���i���Î�/i���a�"�Y����t�*Vv��OR[�V�a�a/}����/��
�t"V��43���8�z^R�E�%�cۮ��}_��;z�}��cI�:q�u�r?;�Ӯgk6��^�< �
=Պ@f���\��ˌ�S��c'p8���gQ�����
g�Dpe���9�U�\^g��k
�L�ѯsJ�"�9�Le%Y�����P]K���(�EE�,enI� ����čM��L���U�Z7���S�9<�E`�Bf:��w<�M��3�舜�&{���YZ�f�U�z!���R��zɞuo��D?u������J�-�
d�`pC�q��WT�!FӇ�Ѳ��z��S�˻���D��<���	�Q�������&1��:�;�h�]�x#�͊�+�gn+�4�<7�g�K�R�`-���Qn��A��F��3�Ɂ��ȵ�p��E��Wj�2�G��˿�"��[e���Q.��`��L%C��ڮpP���t�F�C䒽w&���9�<��}��܇}p�c)F���	X�,���F�2iTz�@}��8��u���~�*�f�5UeᏖ����Y,I23� I�H=�1�ͯ��)��%�.�ΔfYZ2&(}"�;$�Xo_[�������������.���;��s�
R������;��b�89x���GL��X�ܲ%�k��u�:m��%�}��3G�D��,�e��������/R^}�>�ѽ��ł�6WT��%ǾgN�����}�*11�ik�)��&c�@��qt��[f0���G<�ꑰ_��c�����	أ�ď8swT;⠕וsպ�s8$��V�a3�E]=�l�\1/�,��,߄Qs�&2���`�"���y�#�h.�7'���9 ��1��4߱k�a	ؾ���jtҮ���D��7���@�f���@^D�;8�Q)Lw/��r���ѕ���.������p�B���~��TIhy�Z�pʋ��H��� �ϦGT�`�e՟軕&�eo���t� $��jDz5�O�C����<�o:��]��R�	���ǀVQ�`�l|�-x_f��.���3#mB���X��_�n��x�@R�)�a̵A%�)Qa�,�P��c��l��T��n��c-OE���sHQ��)d`rUN��@-j3��Y�r���mȸA���]��@@c3o��+��_O��h�ǂ�iF�ŭNȗɑ��7�F��㧩k�ǎ�Єυ���۩{DY���i?�� �tPS���%M�*�DB��OH˶ff)i������8f�����^hy��1��'\ '�83���<@]Y0���˛w��)��U	iӹ�@
��	�3"nP	����Σ'n,�8�)Y��>��f@�x����"�`\��$�Fe&B�!�����?��Ͽ�[Ie�pNmRb#\�KZD�Ma�	K����(���b�}K �T�w�;�����y��R����}�u�#��Z4���!��⹷r��mL=�Ϛo�d�Hx%���}���/�Щ�J[n1��)���P�����^�J�����Q�W� ��'�����нO\�|Ys7�������Ky2j��b]�Á@���mo���m`O��4&o�&��0nc$Z�T��Y�� Ǵ���3��Z��J$̌�_���m��j[��5q�=�^���Z��[i�	���"��cAgɲ+޹�Ks�l���`+�̊}�((s��+!H��>3Opm�4��G�!��,���Z2Ǐ��9�g�&�↸%�`'�$���:oz��(�+�Ѐ�Q�J�H;��a���<r?����}�~~@�4o�b͕]��O��ﳪ�~9B�5jAOT����

�JPs�.��rA�K�ېӯ����i����������$��D6;+�2�~��l��L�J7�8���ﻵb��d�sk�n�ʒ)qC���b��(�1�&�眷
�t\��v<rʷ�f�7/d>W^��A���gl�>s�!2?g�k���e�Fw2B7S��w$�ш@�"�x���h���[w���|�̧g��I�翦�$��T����
9?��L��g�E	�U2Ň5g��W4�]�,��a{[��+���$���Q��?{�e�gy���ޚ������ؗ��*�G\��o�:Ԣ�|�{%�Ѱ�x�ِx�!�R�1���I��6Wz���!�4�W>����mX�ǃ__��۵��P��D��L�b�
;.�p��/�q9����� ���nk�/H0n�:�F��J�!�	!؉��E��a�<%�H��$hWE�R��C0)F��¼��8�\xa�����$�8���z����R:Pd;���:+�6(l�
S���1=��e���sV���4�Z�[}�sݠh��􂍕�.7��S��������{�ȡ�Xf9����)&P���DNa�
u�p�=�'�ܑVr�p����'|);���Rq���.�gfa�'��@ $nU�F��'V��?@5hR��ޅh��Ċ6��t7�����L�-е���?y�7�dS^K� �!�%A�O垝^�M��G�ę�c��LX~� ���)y'�`�9� Ĳ��;�1[���|SI
�E+�p�᥊��(; b�aΰ+�is1�*6��߂�=��b#�`ѫ'�רc�q\w��� �i�C� Y�L��������"�{M!�n�����|��)��΄r���U��Vv͛�kl�^����V�b���1���F���� "�EC���<%�����t��V��6��fԍ��Mؒ�i�*�\��G�e�ř����j�U3�}�&
Յ�\2;������	|���6�ꉄl�}C���4�HJ��_۔�6�3�	_���S�L��늀.ۻ`m�`C���=��>�rf]8U����iGx��;�W��u5�i�������Vc&�� ��'�[-%�<�}���+�l��U�նn��h,v�̲l���렜�Eހ�e�u���erz����ya���-Nl����l��k_�R��H������2�%�[��3��Ra'�Z��hT3HLP	l���+���ȅ���TQ=IEF*��K�q������,H�&=�hP�e�|~�Ct�W���u�������v��*�Qj�L*��`tmV��I�Z����KP�"_���˵J�eԜ�yZ��{Dq8[Cs��O�T�@R����9����\���F{�����B�z����Ї�
`:Y�wЋ�[��6�,KX��,�ot����Hĺ��ñ�&:�R�/��4(e���y�r�0������Ls,���Ê$�-�icr��b�jzK9��l����P禃�Z�E���k�OW�?$�G��<�`�9}B�Cc��ޥk�EU�v}��C(с��.���N���J�$ �yna{��vJ���:��@�v����=	�ΡV��AG����v�g���he��aa5b���y�غτ9w�V�AgfjL�KS�fG���'����o&&D�Rc؁A%�ŰU�I�%=�W���o*@�e6&��w�Z�6w������mB(f��p��q^�/��ج@@�v�:'X���=^wЫ2��P�3pF��z����g���/�|Hn��
Ԕ�����T5/Q�7{h�M7���uI��.�_����^�e��R�
v��f}���0�����{�Zs6�vwHy�P<!��.d�c����F+Y���tBbl�^�`O�� }$�S��gx )l`eo����&4�盦+,5|{�B�^��e�#ք��&S�w#�y7K��v`6*��n�ӯ=�Zɘ4��o_����iŵx
c]ω�cx�D(��o�h������?�Q�)[?M���蘊� �8�)�;2݉�����qs����K�Tb����X��`��R������'�����	q9�:t?j5u�%G�FU׊X<��;��Z;Z�I��#�h��j
2�ɲ��4�>��u�/Q"�FwZ���;YO�Ui6��/�E0�iŊ�Q�R��;?�p���#��@ÿ�%���(�uRB�8�x���G[�g�tSH_�J���e���|��]S��RX'̇\9����x�	����p+D_��ku玧�lYħH�q�<���k\&�s�m�ߕ��)�6�rJu�ɯ������14�+�Š�E�=�ف�jNN?�b|as����Iy[��M��W�ւ����c�zW!8[n���f�A�:��UOB������jO�]=|*A��k�?P����UX�:��ua�h� �+�.3涆���*9���X��������4 Q��)mI��w���7AhC[��BK��K�逖�;�l*��#�|G�eVŒ�����sW���:r��?)���e�m;�$o*v2ב�1��$$�����-��+R����\��y�ԝ�1O����m�	�6k2^�]�춸��_@�K��[l���v�W	�$�%ֱ��sH.~�n�%��1�vlC@��x�o�w�ϕP@�\����6��+��gU�d��Ќ��p��5s��:�v�e�����<-�8+����js���	�?ٰ���)=y�6h�;@F�H�fo� ?�!_��ƩW�N�t���
<����-��3<l�k;�@�ҦL��p.4�۰��p�i#��1r m H�'k&��x���:��^�N�����֠ +cO�<@"u�4�� @��:0Eyg]�0�@0���aPisc�*�*M�� T��Ҭ����C?��;@�%'ب���Ȃ-�F�q=m�X
<%	�R8�U��8j�)�.�/4�O��<����ʸ� �=�A;���&F|ϿX�6�-	���M6�F]{S�Ud�_��b��C�.�Un)�Zcnq�4��C��z����'�Eù؏�����FIó���@cEi���E�ʷ�XB征��}ʠ�*���"{�z5����̸Z+��Y�Ү�W����r_l�z�;���-�|1#�2�N�	t6b�c������k6s�t���g=h*���D����/l�ݮi���ْ� 3�B���W�=@�ЖHɴ�$�دaSBĭ��[������(�
 �!<�g����Y;�6���gP���Sބ�Bl�Hu�U����b�!G��%�
<�C�8�����Z:�+�+x�D�5x��=���RK�Y��ֿ�Sq��0
���
JoB�D��fZK�зH����8)w8f�j��ϰ���9���3�^o/����qH�$�MY��4�:Jf.t�N2`�0L|���A���v�l���ț�������il���xƏ+C���ǔzs��_���6󞥪��vr٣8iU*v[³�^H��@���4AZZyA�e�B膋�����`�i�\BY�p��*�K�Q��\|<��a��&D���@����$�]CM9Qo��J������V6�%;x�Xΐ����������}����`H��2��i�� �}n&$�Go��C��)����«ƌı�U��׿Y&uXtѻ��g$F�<|U�C�'J?���[//����P�?ʊ�V�o��P[�6���Ie��"�_Ep��y��+�J����Q`���4JUl�����p:��HSqb��2�E�N4��:$D��/I���'ӓUMZ�����v�U�b����|=� �-�+�� ������f�[��L넹p~ <���(����I�Υ�-�[���6pT�#k��hEP8s����v-�"K����5��,�l�$Y\'���c�/�Fm���B�i�FM!����b�M�ۆ9C��VOS2��������$���?y��>�kϭ�en���"�����>���k�BsG��|$0�j@]BK[���3~�yR3� -^0�cs`�O9�i�)8%�j�R�p��
2�9#9����8\�ǺK�P%�	�_�zWTi���$q����S���v�>YZ.B'a��6T<�Ʒ/"��L�y�* ū-,�6e���G�EqBU3�t�����K
�ч��
}�D#TSta�H��C��p���H!8��Q�b�r�p9e�rX?��=	�c�u��T��z�RP�>�v�9b71�wWi�#�[*9�����	n\�(��X
GA�h�c�Ƴl�,�{���[���Y\Q�M���J�&-_�<�<xޟ��D�ˡ�AH-�/6Q���t�|��*�<0�6y��~iS���L5/�w�3�%X�C��⏣�P����ѱ�&#�V�?���n�e,�#x/�/m��S�#�ۄ��`�yFi)M����j��t���rNr:В�D�aͽ.���Eko;�/�Wa�m�E��s;���q�u$�£)�q���6�rugŢ�}��#je��)��|:p�zۇl��g���x�˂�!f��yZML=�� ���
�~�^o#���U�ꪅ��x���h���W���u�A���z�r5�\�L�������dpv���J~�y����c�F��+W�1�8��O���J�OǬ���M�V#q�����\\��d)�<Ѵ�h���ԦTւ}2�-��,�=�/�#aY�B%g�W���1In谙��vA"Ȧ���σOSV�KZ~�եMV��A�Ii� -�P�CX�c�i��1&VO��Hx�O�u�/��g[��,�ML{�Qɭ�̬S�t�!���)�D��F��%�k�uي}p��F��P��-4��r����;�I^k}�;���a�p�$ ]\���n ���x�[ߠ��C':%F����%������p�@UOQU#��%4E�	�),��B�fRSIv�a�\N�/���_�Ly�Xm�]�}��:����&~¿�������h'��\1;��!�f�d��]�*.���r�f���ީ��c[��,`���x"6���c�C=t��G��Ю??	���=�f9��.�RE^���\���20R<W�w^E��x�=�z��A,��?�P��J����  Jb&��Kx�+uj�t}WSEE�:�yc�Y �;��A;�}�T&:ʖ�H_������n��2[��H� {�Ė��3�⃵�9�ܴER��n��9 h�rX��\�G��XJ������黰G��N�5���d��'g.��]�T3̗j�����~X��>_��m��#t��94�]��F��o��bQ5��#���1m3��5D���D�U���ث*�'c5&p�e|����/,���w��=�QT�/W=t����ꔘ/��@r
��GI^�fl|9h/:�*G�!�`��R��EI��K��-�ht�Ҏ3B�ɜw?���}��ͧ)Fap�-���|�~�Q���⛕J���1+c�Cz�6*���EG����)��R��#Fj���2;�8���J��2J��u�m|��s�x�
9G�zs9��o��RXO~W1K�f=���M��O�>('8��1Zz��F�J�;EW�6O�T��$.��X�Ɲܫ����Ύ�,�(�����ٔ��$�e~y��a�!�Z��T��+���[�G%�a,�ж80�=�L��]�|a��&C��K�o��0q7��w<c����)��,ը���|'l�s#��$!�.<T~���Ee�E�J��ӥ��>U�bg@� uM�Q=��6D��oL�s�7;�'?�Q�RH����?�������g�p�
$��뛡|�Y���J�l~j�Z��GÈ��6 �������b�o;���R㻖&z?��v����8QOl�.p���?����HxJyve�?�I�Y��]�!&��R�-��Q��Ғ��qj��*s�ι��*ZP&�E��H�P�����s��6y�r�Q��o�H�U"J��$"���
����3����߶J:���9�~��
Q��[�E��@��K�1j/2O�]�����)�����H������O}�B�ו����v�=���UG9yFm��G`?�e�n����jI���ׁ�����Z���RX�V`���ώv>����P�l|gK�i�qi�)s�*�0�0���*|ÝR�x'��ncX�4�_���a������K��ڜ��4/�8Ĭ�N�!�&IJ19�`J��m��d�+�[��S��I!)3S�g�DNP�d���u��Fޏ�6��jt4���([��ȹQ!�a͏�o,q53�F��[��ۦ�Q�]|�˱
#}s�ȏ(�����q�r��_�TK�;����e?P�	02�� ���/LRۆ�_��j��Q,�v�Z��u��`���C���!̏�(��]F�'�'|*J�E�컰�H�0�W��4CT�d�Ps�P˟[�L~0�0Q���{*mi|�l���q#��TK�g�W�f��<}�*�A�����P�~z� �|A0�^�����j��=��:��jю3ha�̓V�|.�Zy�.V�l�Xw\^����e�c]	�k�^��Q�$�oRزփ�Y�b�R#��l7tR�aJ�VTx��J�ګ�T�G��/8��q̅fg�'�?N.�p�-�5R��J����H���k7�2�8�o��a�4!�����j8�PrS���|�0W|�%_Y��g����I:�4��*����ǜ(���"d��t_��s�V�o�R��gf{I��CΟ��vEr��<�j�qhj�\-\�ԯ��o���NB\���%����0�����B��>���m�o{��X�Ȭ�]����[�R�!�u���m �#wXM�cpȳ�eQ�w�4T��[�Nw�j�{~2�x�����]������S����[W&�n���x��3󺭥:���y�5p1�;��~.)�������4&\VSD�D9M�n��؁�l-�J�gK��Lk��<� �`�u���.�{�AX5�"`W���](� �jU���X�p55Cdc*YA�;>�؊~�}-�+Ǖs�5G w�+G���|b�mG�(�BO>�#])����B����4��6��1�:�v�{k���	���E-����]�1��~���M��J�f�-�D���
Z�7<����6w��)-�I�M���wr��I=_�ͽ�����aw����h=���y,׍�"�e�,��ȖvH�qK��
q6C�N��)�%��&3l�*�/���Z(�rZ��)���}c�N����߆�<�'۔v��T���9Oߵ�V(�wQX�E(2oJ���b4���0�zxt�QI��Bm�%3�/t���k�*��'�)2���͂�w��:�B ����u���޸��9���i1�S�v DvF����|~��7��#���FW����J%؇�B�<lU��ߩ�y#���?�SSw�b�����Q&�rd��LP�~��"��u��c�Ð�)p��E��'Ŗ����ʎz ����~�.yn��+]��>�ۣ(!�G��d£u(�����X���T
jPxvd��
"�%�'�~��]*E�����\��nk@0��u���@���ȇN����3�H��� �WU�n
S�v�'Ȓ��s���c��?k���b{2$��:�|�$��w#9i+hh��7��KK�p,`�b�}UB̫di�k����=F˦��׫����v#�$�ŏQ@��9�yE��l�;w�+�B-o^K�.f�P�K��<��S����=�PJ�UMc��z�-�K
c�L��uƋC-��:���`i�����:�z�M�������e�"X�c��^��1���r�h���`���냇,K\�& ����}aS���5:�-e��Kh�����k�O���<����s1�J�L. �ڏ-�n/����ٱ*-��-k2��&6��_A��,o�����zA�W����Zԃ�����@�\֑,���זQ���ᷕ�o�7d����K�ݦ�Mq6��jw7(�@�y�R��Y<�Jeᢴ뀢��W��%V����H�|��I6��w˃:#!�㮭p�0�H���Q��h	�������	S��h��)�����j�0(�
kR����l��6���
L� �c��2'�:�C6��į¾OD� 8�m���Ed�G����r=#C����X�g�l���`i�g�hy1���p��э���b6l@��<�>s3_�������m�G�n����̻#�1?���fĝ)q��g�.�DD��%�JK��ޑ[3ٿ�C�� }�\U�Q���V��&���"�iW�1�j�G��0�h�U�����jd�L0흔,���D���["[���aHe��&��A���n�u����e^��R8��j�����G��s����P�uUR�"�����W�E��P�����K���Bߠ[ơ��!����?m�r�P�o�e��A>�ѲZ	BD�/�*��M��` �7ۏR���P�$�G˶D� n�mJI��r�LHُnr�������������vߤ�JӃ#���1�^C?|B�?�"�*����K݆����D�9������kg��cq]z4ЍyV�}l#��l�}� �����Zɐ��2�i�o�	�y��\A�O���3����:f��o�B�#��z�~ ��s�sޱ��<��au=���E�Ml)k4�/�Ѣ��VÒ�p�`�*�2��Yt���4�'���6]�0#����#��.#��Y2�_��
C����t|?M]i�z�wB]�h�⚀�O�{E{&�$r�0��g��ƴ�Ġ�#�7�4��o�����.���h!��;�A�_�J���=�Y�;ʥ�{��4X20�B��Y(wecn�^���|Ȋ#�^�H)�b��w���^:i*�}������rc� r�H\�(���H���6ib[�U��;I��ئ)Y[d`��Ցr�� 6�*�*G]ŀ����T*��6D��^�7�h�m 	��s�q���V�2]מ��d�8:Oߴ����|}4Z;���9�q`+}@p�_�!cdWO���OA�2�ɩ�s��B���a��^�7�l0��B��i���B��`z���^��恝��~�V^i�%��V���XT�4l�|����`�e[h������e?�W�Q>F6L���PoQ�j8`��k]v�Γ�W)�s:��Z�"k��žN]cm*C��y���)�(��:��e����Y���6��'��o�%�ü�F��"��3�3�u[��]�3���V�ҁI
���$���*�2�0�U�P4C�u��`|��8B��F��͚�`�!��9^Ҹ��b��iʞ`Z{�5�� �p��{�u��kp�����RTn�_��CZ�s�г(ި�� ���D�?Ⱥ7��R.F���
�H��DՂsy��ħk�Ս��9�(����8-�!25G�ѡ~f��5|Ad��*�K��]���5�Nc��^U�ڛ��0XtJ�1�'�y����Z0�7�[o(���0����_���R�GP����jo�E=^��,@�%$Bx��L+�)VC�L-o	�cຆ���i����h�UO$�T!�����k��AjY���ڝ_X&K�w��9aJͰ�����.��\~�p�������;a�&!��IO�OAߓ��w,��&VUgv�łsp�м�9��`F�b��������=|���U�v��qy{-�
�p���[��Ձ���d�Kz��ֳ͉����UP���&!��2������������v.m�ӗ��Ò;cgQ�B�=le��Xda����D�gI��o��Ú��f�fc/�-��^k.���C��Ș2
e����������>��(r���)z�'V+5�mgʳG[K��2�|3tkx7�2�����H���@�T�v����O��с��:��r���|!^S�;$���&戦�ff� ���cS$4ux�MX�U�ۼ'�B��_`�6�NKF��~p;м�F����TQ�gw���������P�ik`4�,�À#ڼ�^�<�Oϐ ��՗�4��}������Q���t+����³�:�A�k�[M`j-%��qٱ̚FɁޣ�k�L�z���4lL�{��8׼y{��4�k�$���#O�%�W�!g�1m�b��fؿ.�o��M&z�ˮe���7)�)li��n{�]'.�a�쯇Op�A�{!��ɪ8.J=+���6����=W=��>��=y�;���H��ʗ��I�B[��ƸA��[�"k�%[����������V��~	�	=VgG�Ήţ	�|��:e!'}5�U&TC�����suZ+��x��]TN��ǭ�E���H�{��p�@�	$�ή�_9�0z����3��N�����4����+��ar���Kfl�j��g�	�X&�|ߵ8���VOEʚ>���nLE�2TMW��* �Y7#�V=�,���=����ҝz�s�4�o��wO�Qs��}6�ZË�[R����I!p<kc��2���H)O�b(}%��ݣ��-�u�$�iF-���*�R�:r�v!�A<J2G���e��z���V���̰��A�e@��l�� ���E���h�WI�"�e�w�=�??hi��NC:�'�^_Eb����x{~�"KK�=���ԧJ�ĜP����얇4F��.�K�77[$�UQa6�xx�Wk�2*��&'�t�Mz�>%�*�Jf�(��U���7[ .�����|�Ԁ�%�]�tB����P׋fiIt��Ëa�r��V	����щ�?;���C�dpf�h��gbNgu���f�I��9��s��� ˞;��z�Q< ^���B��5<4���7�˯��U��x؜�j�d���9fLГ>'6ctw� m�Ѭ]�L1*�m��9f8k�~l����#�вq����#I:�V:�TuT��v����(o��Ӷ��k�{�IՖ���o	��*�Uvo���^��#�9���z�>�_g���~K�8d�w�z�� ��k�xp�L-w�O�4���!�Jλ,��x�[b��%��Vh'L�d6�?���"�<w���6+��9�����J�1�tq��I�c|4ϡ�iI�>��W����aha��J/ցSom5����r�4jk����&%	�K�7e���e|�nv3�W��Zl>��aY1'
�ӎ�޴Y���Q*)��]	���|[�����58�{���ܭ���Ć���B���;A����E�&`��6�u�W?"l���ZJ�a��e�P\q,��A�+З��8�Ai҂|��l ���E������r�4�X�<�n	��ؒ���[<�Ǧ�d��B�G���t�^W�oQ8̾q���MQ=��u��[�1�S��:=L���k=*��� Zצb���ֈ�ayD������m��G&�άz�c��JAo��hUvt�[����v�L j���f� ���ޘ�nش�<�&M�l@�O�ԖH'���ǣD���XMIYս3�QX�}Z9|L't�aJ㻻��{ܸJv�߆����A���M�!H ��n�Z�D뒗���@*��[3ݚ�>�ŉ�a�ǔ�B8��(�u|��l��:�E�k����ܘ� �^�T�#s�z?�\R��c�Ґ[}���6�*�f����e��=i}Ct\�8d?�$�f�=��&,G��('��AqY�"�h�)-Q�V���5�:K?����eۜ�'ۚR�dt�!X]��������1�П�nvf�Z�^��:�!�-K���{���JFYS�,�18�(�;N8�1M�C�c
l|C	#,g�����G�/s���g\�T��"��,� �S��H��K]hzo����ěP��T�%��HGF�T��-���ء��,;��%��P���X2^,��)�pd�Un�\�j���j���\��\���Zj%q�4��x�� �Qg�,p��F�n�]�G��ͨB^n�쀧��qCZx�{TŐ�_�����D~ߞ�e$E%�(c%��	B�7,9��z���B&�7Vҵ4�VH0��Ss�+A�zo,�c��7Ygh��|u�$}��	�6�ꕯ,.g���q��N7�O���.���I�KRrC�H{6Kwmŕ��RT5>�vv�����2f����{�6�1�*F�M�l�GL��#�u���rhE���p*R���=v>�(rN)��mv���8�H`�%2t#X$�<�~��@�DA���R�ڰW�
�'�L�o���r���<ʪ�GA��^���S����+��I�*�ܡ+��F����ǬH�Ȏ� �GM3qbx��ʷ�����vi\/�� �%������|��PݘYj���*8Z=S�h�n��괷o�[*���1쏧�Z���^JGI	��Z���'8�6���EoE�'�<P@U�>D�AERNR� ���a��?H�S��F���l�t)s���>
'������CX�,���_�u���ɇ����ŋ�;+f��K��\H)�;8���s�7�j�~��Q�=�BW	�d��5�����4��h�Ķ,R�S��d�6���fA�Pށ�P������\��慹U�0j4�A�n
-���C�
�8�%�������ne����B��0�X�9o�{1�P�,.^P����W�@G�>��c3�)U�G./|�����3�DU��qn�7�YQ/��{+��	�X�O� �ʔl7��AtV��Y.kcL1)X�Aň��\��=�NH9�V��<�z�
vO@`�L����3S�L�����ŏ�L���W��hZ�g*% 1q�甑���U�r��Ƕ��r�u_�r�V��ǹ�-�|]1Mbf
��c81��֜��~!aŋ��G�ȥ���e�]�kd� ��g�$we�_�!ԺS0\'_
1��+)>�N`�r�y�P�1��/X�ߎ*�>�^�x��#r�;�{�#��X���,ZnO� � ͊��r�/k�sN��F����n ��T�2��[�QA}�ȥ�?�No�O�$� ��x�א������A/}�:�M�^G�!��zw0 ~%TK�Pk�Ry��.�3�$r�ņ!ယ�8�4Gǻ��X�@/�/L�y�Z�
�h7����ڞ�Wsrn���5'X�9���vԦn�h!�����&���5��]m�A�uS#��Q�W�� �?t���7˧�Ń���s��f�����ܤ<$)�wqJ/��}{�Y.%�&��X���ΰ׶ڲ{-3N�[v��FJ�ON���)��hUSP/$/�f��_��B����ݦP>�T�M� Tk@�!�}Y�+�+#�.��o��|�I9 1���j�:b��w�D���b	l	Q4��;��6phj0��^�%�����W��̺�XJ��Q�0m	��K���b�^d��
U@XQ��=�Wð�xc�Q3a�:HH���DS	[i-��B:�ܿh��A�6�����#jlU�k�{����%�2��4��J���F��x�g���j�����P2YV�J�MQ�Pg�]v��NYĵ��L���vX��|��UASXVK k Z�ެ�C��ǳ���L#�ᔜ�2�>wU2e*m�7PLz2����ϸ�M���Kw<���F���CQr(�%�7� G�a8���ڈk��H#X0�	 J�?u(3I���
� �
��l~�;����[X!���6. J�'��צ�C��Vn�S��Y����*R
�2�u�=�za:,��F��ܯΗ�m�砑�FhsO�U��;u���3I��T�ilZ�HYY�MCM��_�5�P�y2b'�ر�*�o�ʍ$�Pq* �r�DM�b��im`ІJ��6��ب�%�ر��r���Q���n��2��g�#������� ���umV�蚻��`[6/������
<�ڌ}�3΁B�Xz��8����9�m���qL��ilЗ{l�p��E��@+V�C_���Z>��#���S������U���Q�s��X���d��A>�9(��4t/3!�w�;M�=�.<��mM �[z�Z�x�8���jf-z����e+co-..$#o�B���Nl���K��>�0neI2��4��j���1'<��=@���_�Y4�.�w���������@-�@~�weKP;�b��>O���<��?qT̕U�J��7ꎙ�DglUKࣦ5��D	^�Mt8��,�7=t�Emh.�7�����k;�c���t�ǿƥ-�	)�d��~��&}e�y.�D��4��	�.�ʢ�u�1��Ld��|���PAs��a�r0���eۊ���2����I�n^�.�pV��.o!�U�E�vi�m~��c�eks��\,��[/��ܫ�K1��X�=�/d�-!��G�����{Cxm+b��P���֐��/ф���N^Qf�`Q+_��J��λ�렘����� | �k�D��>��>��s���У����YV�r�J���,ͳi�ʳV���&XI>x��ajNP~�U�)!�c3n��K�܎�q����Wq'���I!���ں���i�wXs�gV��tc ټ�`5m�yD�nS��3���~�t��Q���(
(�4��[�����f���fi�1�M>y쒘(�ӳ�_�B������-���;�!��~?1�'ټ�w�@LB����3�JbG�mV|$(��vbG�'1�����
'���x�"$��]򘪟8��Ȝ�ߢh�����ӊ�'���qw��d����7xry?� ܫ��
�Y�L G �?l�G�<(�ĪX6��6epЫ��5���V�m�?�ta�wV�B�f�|�xx���Ӡ��s�8�\e�9A�1R'f�c�����"����z?q�*"������r��ۿ��Tt�iVtd�#�"�������z@��S�K��J
�B�\jY4��d����&�����rO��Z�A\X�1������ �i�O� ����sA����gط�JDo�y�u,\���N���/����{%�%r|�����k���N�F��lM@���d.`��{U�9l�!�����(XG��7��4�klN_+�b���2��M4��|�H��쨔y��,o~�Ƿ	+3ݙ�X��L�!AQ)�A��[���u�A'D@T][���u���zJ�D��U@��|���Ǒ�'��%���mq����,����Ꝏ,b��T(���rlX[��E�x4��]G��c\1��3R3��]�T:��˅DLJ}�%w�s�V]�1�$�nC�U"�������p�����By���jdsE�ϱ�4�]��^x؎����e�n��W
v�y�ДL=��	=�ǵFǨ�cѼ[��m���d3v�
�bg��N��tk7#7u�ɀ�0|��f�E�^B6Ѻ��"�{y���}[�l
������ɤy���q�%�;]H2p��O��7����~�@m�lF7Ԋbeɦ
7���]Փ��Ӟy���Y�exr�W���*T'��,T���݁���|g���,q��S~����n,Z�lOl��3L[�)��8"{��ڂ��b&^;^��p#��Aq�_�}�]%݋�m���*	GL�>�b�45%h'�i ����B s�.��`���c�hSX����+�N�%��*t�mkb�W�
OQ^�N"���d�b�F4���M�z�X�2����F�䅋ф�\a��ҧ �-V?rk�;�ߋ��X<�������(gD`���2�׻d}�e?��/dt?˵��/[�Jm���peJ��+��όڊg�Q��E� Ds)A�¿љ$L��Ry�J��m�m
?��{����F��3k�:�ʚVݶ�P���w�e���@�W��=QRPT�h�Q�\�}B��8Ly�Q�"4�Ȝ���s>���̚��:S���N�)�S��̒\���TW��T���xC�Ktq?=z�O��Q<xVBB^	���b4��x3<�<�gT���p�m�	��uǼ�~�?�L>8�r4��Sa��:3�@U�䥚�CYes����!���$���$. ]�!�0ώĸ�"JG
�p�ކ����~a�e�b�K1b��%p���b$�u�X�Avi�*��&��u���jf�L���䍫���Mj2��):�^�|^yR�V�I�4�V$A6б���i�]X�Y�;�j��hu1Ld�J�b�CuuN�f��cHG�C1�� ��r���T�M�i𐸤B��lp�	:��l�2-10nxV�Q�;�i��pХ��d�MV@�2�jq��������,�"��ܭ#������yٲ�BoM�/�\����b n{F7@r+���泛�W&4��X�S�7]���"��L۹|T�����e!�9���0�6����H !� !�3���!�ª�SU��������ǲ���oj�Rbu,�����4SQ��jϩ�����0�'{���`��BB����I� ��z�R���lQ��<�
y+23��/�q�r2�S��g2�&!�dR���#�.�SE�$��hP:�8��xE�+� �ˀ�g�H�Bd�q�e�aY�B6���t,��ğ�ޣa�����(o^�E�N��#��]����b��m(ul�{&��J#B��7]����k=z|�qeY^���#�]t�;#���M�~䱆�_ڞ𬒦����=�y>��s�[!��p-Ν>�-�G�4fZ�:�)����<����Ç���?vj�h�Ry����S�6���p��,��p�]� ��7�3[o-%�h_ZEp��9k�z��K��0s�dI�O�)�el*t����uYQ�㣌��pJ���0_��k^�&�P��O������t;��er�I��g����Ւ ѿ�.*zI���f����A')���6HήbQڋ�V�/���sA��I�E�`~n����;>����r(����^_?X�T{��7^�����cT�8�ɑ�8���}w��(�-Fjn�jp��WqL��l�N[�M�7
Fŗ	皵<��1bJ���<hU�~Kh���>[~�"���@z77}ò�njAM~n}�hԻ���f�rkM��\M/��$J�������峹�6��{/�
���#�,����L'#���=qL�z���vU3�"��0��W�y1a�(.�l@�؅�[Gh�։߸^�Tһ�2cD�����ϑJ�O�T�PPY1����7Ov)��&��wA�w��h)uPh�t5έ����
�ˆ� �CLW�����g��5*(����2���.n�������C@I�N�yd��jng
�o�G����'�ԜQԧG:��.<�}���m@�� �������"]��z���>�x��-� �*��@��J.=А4��H_Hu[4�o���%���R�j���^�&Ww��ndQ����gn-�D�B3R{��0#���eA[�Ï�t���]v�3���eJ,�G'j8NT�`�^}��9�!u�Ű�%!���]z@�ys7�|�93?�L14��U>�?����:�����f�f+�4�s���q5V�m�����O�m0�2Ҍ��w�v��Q�hI�S	y�E�7����[n5	{y�����粗F^�J�B4�l��BX�o��L���,7u|�diLB���	bs�d����Q��a<p��Y��̓f��&���]��Fk p��Vr,���1����E��b@�4�_��A��	�B���J�͚�se��1²���Oa�c5�u~4�������T���_oe��m��R �`W�%o�������y����oZ�{B�@�]qBj�hOpx0��:{h,�[0~��sO�^�������i�I7k�T��Z�IO�h��gd�qz�R4�ai�C0���o~q�����{2i[��43�
����m�� ��(�����֠l��-_�!res���& �tų�_�2��{Z&�+���
�r������@�yT^	Q���B�Rp���,�|L�8�Eok:PL��>��w��'(mС&��g>Pi���t�mp�S�M��˺�k��u���8)g;;��NքQ�P S����hMa=x��Vr�d����}�^Z׷�u��V��v�%$C�^3~���zS��OVo��Щ�r���씧�i�0n�<^�.S�N=K�_"�j,핝L�i��Y#wTx�PH8*���Y|I#Dsºx��BM�=}��c�)�r�:�Ve�\a�m��d8����i�C��t+o�^%ˉ݁Q<<ޜ[�4�t�xĩI/h.-u�&���N^�)�����]5�^��Y�Wײ���k'�!e둂^uA�:���4`�{�������@�"Ƙ`U;Ͷ"J�Ѧ5�!՟�&$��j@wr��Z��`,6�UL�/����MC/q1�V(����j��:����Q�20��r!4��(}-IO� ��X�sy��L�V�f/]v��;���f��O���-�.��"z��cפ>�U)���G'��٥�W�Ƕ;���p��q��w�d�q�$���JRP���\�[����'���^���[PKR��d��Ty�m� lh�l�	�_+t|y�w9�3�:W����ԗ$GӞ��;���O���9!R�9Wm�XFR�����ݭ\|	�.��1^�O�
�j��!Y�7m%�C5��U`������[z��_7�c*3��������g������tD$β��`n����6�1�Y���X=<+�!�r+&.t
2%��kz$=��I�"��bYm̸81����r�pT��i��D!@��̎q䕄L�Pf�!FI//��_��)�6x��5XDK�5$3���i��n� B����,b����{��t�؅���f\?�Y���7������SK_=S���]r#xi7<�DF�~�fm��7
�>_:դZ��B4X&�dR�C�Dk�ɖI�P����p�f`7��]f�?��Mu@X�G��y�M�A��L��A��@tJ~3_M7t	�'~cK��:1�9�k���|@�I3�n9���K�4Iフk:ODO%�c��|���p��}(�"��"�N� Lq��]�L
���Oy)#���W��`�Y�jbΔ� Ё.w �����.�9�(^<�-Bȑ��ư6b��EMW�����\,K��֚�d��#	�1]OP>Bɩw��4@ӴA튩���)�'<�9��ٿ�Н�I*���_-s,ɍS���[>�}�6�Dd�Byk{��v��`�~~��k0�T��U�wS��~��2*v��T�j;=?�w�<��'�2~e�;ev6�7k���y����1��lin���,���!:M��������cVC��hT=Y��7 ��rC>�{Cڦa�ԛDhLrw�}�ޟn�s���f�Ef�x�HR]��T�����!���ulV���Yᔫ&���Ԧc�l>ʚ�������&���0d��ۿ�q�jh�\ U��l�Yn��X<-E|�$�aS ���A��K�,G0+����5����U��ME�I��(A8A�A�;�I$B�Yn��R�A�� p�Iѩ���@V�6��DF��L>$���QԦ�Y��\�K�8 �RO�����C2��]�/�@�yx���Yq�0���k�L�����~`�<�q�jz���2;�����s��[7V�Q	|�!J�Di`jJ���L3����h��{7k��aöA��O���[�,�&��}�3���b5c�hY��P�0�����j0�塈@A쀡�Ц�5 �#����V���t�ȽE�H�5�:a�l�)��f��̱�˧��L$��?�3�mO��ڌ��Y�?�O�Ӂٽ�$�Z�.��kg	w�멹�����1+!##�4�ؖ�v��?�Rh7�"
��(H����%�)� �/]�Jlz�����q~�WD�W-Tp�M�у���gy��U�ܼ�Ɇ�؆贋F���de���	����wms���J��!>����	8챖޿U��;�D ,k<A&
�$�5�����Xm�_\s5��^��j��SW��֨���U��z�l�1u�gQ�ª ���\z������K�q�K����da��_��-����P[o��E�t��Y:����t,���r����g���\�`b�2�7|н�q[��A-o���D�U	;�v���Ђ��x�����i���f���i���$-�N���J\^�w#���k���t��o���-�6�/a0i}nHB������������/Z b��Do�T+��V_�K�S�e�O�o���9C�K���d	�[�F��?8�7=�@n�s��$(#s�����Pk�4��Q��<�$�|��%��J0�čA�;|�ؼ �ӫ_�O��f��]��l [�qWc��m����ן��%S�K�=����^	c��l����(�����:$��n��֚Vm+�/ͮ�Ju� �_�^�ͰV��v�_Zfa*��u�4��};>������@�KIl2:�L2ǂwe��L͂�F�X5��B~�|�4K�&ܼ�5@�{K�YI��"�^I���&��vx��h�Aj���	�}Us�6���m� �����&��V /����R���uu�*�_{L���7E~H��W=��S��l�Ա?�4a�C��?n�9���X�����!��Z �Y�&Xֽ���s��t+���DXfГ��q��	߈�� �5O}[��}v�4��lRr	�:�E��nk����=��ZO�L��#��[Aoue7ϔg3��֮+�z2@��5kd���w7��҅6' g�Q&&*!��^.U:	K�Ȫ;�7�O��Ю�Va�j"���Y0���o�i�m���u�����ĕZN��c�6?X��Hw�v�S��Z�(��A^&�hSY���>��G	��N����Da�?	Ʈ
�''��h|���'x�M�8{S���
��h�'�jhS_4�­j*�12Ci��`�]J�*���Sx�B�{s��.uP�n���T��6�-o�ŝ�M<�Q�ge-ˠ�<�@_{�'�B��8����X��V�q&�\I�z-4�Q�ibDL}��f�z>�v����S��2"��#�ϼPj�p��h&��K6�XZ��8ߪ5�?�{�$�q��m��{�"M��s�?�k�E�W���9�M�z�<�w�Gz�<������s�N���@ᾶ[��4'k�O���
=�k�U<"�iuM�-�zr�4fyQ�(_�ĥD����˗�iX��U]�v�5T��7LX&4�8\�é����m����,�e ��B�*�
8��ho��g;�-8����ߴRT}��� 	������o�tVT�(���0m���(^�(�Ύ��1B��[��̌+����zZ��H斻��Δ�*a�8h�Z@�ϾI{���H��ς��w���K�m~DQN���\ \���2W�M�B�ۛ������	�����9�0ɼ6h} �f��V�µ($z�v����Q�ǾC�!�x���Q����0 a�5�-���:Ѥ�t���ڞ�&L��&��m� ��3(;m�gh�
�I����y��*�oY�� Ҍa��s�;>AV�����_����@���<|P���1"��cF���(�L�[�-#�v�k�g^m?i�a���
�YV�c�q\�j�B'��p�ϫ�ZD�`�"�f����\r�v}kq�5�`4��9MM�f�yR�l}���q*DI��U���׍�<�/;��4��/�	J�v�R��B�ݘe�RE��� *hxDjᵡ99/�4aצǆ?�-�Sˊ��g-W�6s1�|&�y�Û����'�^�G�~�Q\�8dhy+�*�!��x��� ���	��cN=dn�if�7�Zf��,Q�a�m�@4���*bԧY����re.��s��
� ��5�y�dʛS�<	��^�+�(4��YLRf�8�}�4<����w����2ӯ��M�H�,�fݮtj�O�q7�m+��jI.�p��ڤW�:��g��6 C�L��E��[��
gTvs:\W��ﮭ\�<�8�����嘼w؋�}�Y{�v���d�GHMj;�!�������n�9���V�2aԽ[,�ے��C��4�$�9ظT��C��k9_X�X����X�szxiNB�!S�09�o{�5��.�����vyG"pm�#���!�XAW{�WΙ�`��;[��r��g↚u��
\��Mm�El�,�|�i77��^��}�64�B}V�F��<��oQ�=<�x�+�@4�<�f���ՙt��%$O���UI��4lȂ�_Z:�P����]M���B��Nk�� �°�|\�\-��t�e(";q�q�M oO(�bCxe�-���r�����WL�&�=Zezq����IT㪪�)	�i�'�}�X����+�<�����K+�	�_T�������H/y��.���y�\@�o��G���HԅY� .�z�?*��@�-��z?a�U�0�=���� �W|L�Wg}��O�Jų��l_�r�&ͨ] ���)�����)����-?k���l?ƛ��Ȁ�n��U��G��^��eF�N���0$h�r-�Ð!'�ӺW����� H���m�:��W�D�2�ET��6 �V��zw��Ez�ej�����G�'J��&�{�����z��N����W�,�#��+������B����Q�b�v6�:���ߧ��Ս�Hm'���8*�h�&@�yMQ���RÏ����z�>z� �^�
7�h�'�&��kq����/V�b8�Y���iD�{X��L�C�x�5Ω�Lnݛ�ާ�E����,&#���Pf|33Ց��a�g3���J00�=�*����ZSY�p��m�C"i
��}$kwn�{d)�BgC��ԣ�25|/���t��`���Nd�2�$�7�掠3\|�6��̲� ��b�|�m�3��-� �R1S'�Br�L����B�qi�7<5~��,�zV7�����ө��my�U]���K��$[x+��qp����`w���qmt~�1��`�������_��41#������Ja.b�}a�i��>�q6��� �T�O�jE�v|1:�RB��{t��nFXF����1��A̈)�Wdu?,�<�I�5�����by�u<�6Ɲ#R��E� ����2}�f5Z��J?����,_�R���������:9��ŦAW��z��ɘ~s��=�(�".!��tq�V�-��mu�J��x���,���@�Ή��KJd/i04�⃏��S\+�ң]�ZE���!.���![��@�X���G�X��5-eNY��𒄻"%�	���i�&�<|cx袗��U�X&�<>��
�?����y�zz����̋oH��(��g����%d4���kR�;�G�~=���v@mvK�@g���t�( v�J��ץG�xܤ1�����4q�~��3W*�d��W1uB�d�f0�C��x�㪈��ω��$M�~�M�@�M�:��̕�wc���Pj�i��_VI$��3��-�9��Y�d�% V��緿a���kI�,�������&�b�y���>��e��� ���[�z�����!Q�i�����[գ�IG�r��.t�VfP��Z�����N�N2�8�/h��i�(�������;?2>�<��;��)������%Z"��7��tk�hIf@�:d�~S�W�{������8ߡ)D��o}�.�୍p�� ��D�m2�;��)�1ɚ80Ӂ��r�8����ՍY��!�ɪ��n��%.�<ZT�s�S�\?S�_V�Y5(Z����gԲ��:B2�tou�q����v���W��zs!:�e�![m�R+�����7�Y��Ԙ5Rm�E����D�n�>�� �'~�)�T��M2h�`�A�^�y�;�vz�&�
;���t;s�<c�RW��H6Q�?W[��J�e�r��'����������!��in�0J�@*/��Z�s��}�w�2�W)���Yy�%�[�Ţy�F��>�Ƅ�F7GRu�V:�Ͽ�����G���v�2,�Jue�w׃�}g��?��ت�D�Fn���ʣ"姷Dp>�3����H�}�A��Y���Z�Tn6j�`֥�d^9���@�q/��;���sр��/X�b�\�m�g��8z(R��ڴ��$M 1lr�l4omQ�ܵ����^dUf�lH�π�w�j;�
�H-F6�X�l5\�Yǉ��G\�5!��� @\u�������������~�#vMUa'�Pn��q����Z�$0��=o��Py�U��hƲ9�����p̕/��)���@���c�я��CX#~����?F��u3�ڡ���UX�m�>F���
�|��6a�G/�*���y�G;U�d6hf�6�6�7Д�T����ĩ����b��\�
���:�Q��>��pǳD����_����xjz�!�+�c�'�~(W�]{�E����[���P���\��+	C�鈚��M�ikc�,��v��qoWmf�F�f(���s뛔m�/��k���1c�̭��M�'�P��.?bpaO��h.��4�ь�1��p�%�d�@�2��iˣ�����)9D�UΖ�K��e���)��τک�|Nߦ O%6H�Y�7����1O�~k�o��jɽ"���5mT�x�u�LA��6j��t~�[��H �X�$��cжb��%�Z����m�)�������-J�^`��(2�+	�D�v�RDO$�F�vq?KN���-�ܡ��J/�KY����	�A:��-��a��f��DJ�b�.��+��|l{�V-��<�=
��mR6�����+�]�nb��� �A�`o�o��W��'6��U�l.g RX|N��<�+�o;�?��R�!����O� ��8����9{ ��(�%�2�G9M���K��0����8����Ӝ���\\=�>ge�8$y	�ځ���/�=�i@uDĥ��W�c�nTc���.���	Pѯ�b�D�*+���kƑ��♪����q�h�$�)B`���0B���q����[q�6�@-���T���H�݋�K���3c�)�����j����i�6 i�E� '2_��L��a���^CP�'ik����'E��2v5D�ġ</�l�l���i�o.�w���'�[-�� u'�S��_Ϫ�\q���+��7a{�1'���My�V��ʘ�ǭ$�E(���;CPf�����{�w<����l8����!��7Mt"�y��y�=�m�
��~�n7jioQ�
n��3�,9|������D�V��]�T�����7yع��ک��H�z�Y:M���6�!c������"�=�f��x��Iy���n� |��pKŎ(��%��eg����M�����{+�+��G?���SoWtz�p���5Q������>2�(��ps*�ϣ,�,���6��nu��O-�iH�D�zݽ*�dA���ZS�l�hd��w(+.HStK~  Xnҩd�@��3'�F1�i��:bP\&>{�:�P�ڮ�?����lC��IK-5`��2`�4M��f}�\y�|9C�A�蜆�[A��!v&>�0�w\�we�}C�%a��A�Ґ"?�����Cns۱�6��ޓ����&�����2��;�F�H�uڶ�/�u�R��7ɏ�C��[V�΃i�����G���khf�5�:ט+���h�ӊ�%�`�
�?%��x ",+�ܠ�ĬlDy}�:�tǲ ��~2d;|�<���7��N����DhX��o�'l��GԤf��N�0�5���ߧ�_/�7�wx0�|��sc��IX�q"��Z�Y�u�tV�GW 2~�[�V�;���vqІ����TS��'kh�9Z����v���w"��'!����
��|NVx��k��l���T����iۊ�����I"�R@�=yI2.�1&?����,�X�.o��	��fa�N�j�u����X~���O�8X��/�<y]M�SƄ~�.��ÿ
]����A-N�N�Xjm�ܐ�c�֣U�i�����e s6�t+��~��x.oU�kG�����@��1���`'�f/A��j���������)���bx��[��H,LᕃvS���K����/+����'��ç>fb&����R�(�j����HVAq�x"�����x�,󰰩R'R:#[X��Y��v��.NN�Wn������:�1#���N�'.mK�<�a��k\�}�F���e�Bb^�&Um�J��/CQj'�ϬE
,�[c��T��/��|��,���ˣj�>���1��⪰�@n㞷ր_QH��U�s\�m���ң�@;���'e����	����/�F3[���2md{��-`܍|�����@o���{<�Y�����JAա�7�S)�d��:���]�Juҥ����(��yxX�B���_ξ���	P��z�P?v"�{r�M�>�k0AZ�[�59$����n�r�-�?�d�\+3�Z���ݿ+�/�F'�2`����������n#nvU�a"��eqj�\]����pj?��%A��_	猖����<�z�}#�ɐ�[�p*S��pu�,�c cc���ғ��2�<�����-iIW���%��w<�?G������/�/���j��l�
�5��f�#m�T<��UC������?�sU���]jJ��V9�&4�UI�;����%Z��8g�R��>'R������ϝ�h�,dۇ��*�]($�-8p��1����~�JV�� �ӎ_Q��J�!�
����#�O�M*2Vg��'�PF6�������4�DPn�ޚP�D��@�@]r&���M���y���W��Q�_e�݌�w��[�������4J��g��)u�:2MT��	4K.sBzMkѠ6��Ņ`1�Z�����y�����Efyh����<��9֔�V���.̷�Z�|�����L2��5=���v�0�b��ė\�Q�IXr���ԥ�ƃ�=�����"C��kC�&��>H5ف�ŨZ��H!TR�ͯ�k����Y�-�'3ٖ�N�꿩����{9I�h�\�����yӱ1i�pΌܛ���w��܋`�Ju?�w�~��Y3����1�)�����ҽwuĬFOT��C�"|{(/�PZ�d{s¾'{ԟ�_�ȁ�gM"�j,���5�����Fs���S<�v�r�ӱ+�%E����j�d갿F��$[ٯ\�I(�'��v)��`�BPL�ǌ��ħ$�la�:~q�#/v%����i)B}�m繷S���Cki�:�����cfR�ǧw�v���ߐ����Á�AX�zIb���X�Le�H���J�s��;oҟ|��I�e�.4;�\Y��t]w��#Gj{�((��*��e=��B��r�<5��({���U�7�u��D��]Q��Mu�y��G^��B��	�[��38��<�*A�gT�qY13<�ꦞj�a���P�u�����0yL>V7!�D��4������aS+�f��aŋ�*�'\+Y'�v�W��# @8r���F��#c�Q�x�P�wS��S�RY�	�2.8��,t�2q��[Ů!v�����"y�|Ǯ�8�=L�Ꮝ��t�@�<B�m�g�u��'[_�@�C�y����1d ��L"��m��Ԛ˗�h	�h�@���{���H��
�'��)K�Tp�,�:��5���G΁=bt�d.��D�Gr�����NRGBYĺڱ�ba$�"S���d�F��Y�l]�W	v�E�WS�!��n2���]�ǶxM����M�m:J����Ϧ�"��~�F_������������s1��wv��)�/d4M߁( 6SO�&�j��[�0u��(��l���۵����#��>�т�D�(�!w�]��I$4R�'�(�(�L���e�I>�(=�������K7g�2}:佒K�s�@F���&�r�ޙ��'B`��_�����I�O���<�7��T�d��{���q�St ���<��?��zE}���wdX�@�U��_���^N�J 2��&�|tLx&|9�z��i��VL;�C�H�8M#R��r,k��!͊?��DawY�{��Y �2�s���_�s��Z�D=�T{HE�M��-?�á�`c4&�Cu������qQ�r�f_�D�օ�p@�dI�q��z�[��FȊ_"%wo������( �>oM���E�鯶!Pc�/nn���s�o'߰/�l�Tb_jK�;4�l�;�"���%�x0�<[X�UGSE<��1�]$�Z
�m�]2.����N��e��o� 瘔{�����NC~���M������mg왪���+q@����'L@�� �7���2p�.x?��6&��,���1�)S���A��(�Hw��PN5�&��~
P8�~�PH!���X�y�z�p�H6�G�����U��-fA��/JA���7C����;'mM-WS���P�_�`�@���+�`�x��y,rV�) HF�v���x�q�=8Y����B���W�5�����'����括��򕬽J�qM��0�0�7�mX�G�q�N@�e������Oe��+@���@�B��,%fz7�%�T���$v�Xꄹ'~��gXo�m�_�!CD�XHBoc��&����:U���F�(5�,��j|�F6K{����u�m���\�\ĺT�{Q5��� ��mfv�����l�gZ�K�>��;A�/lG�oi����g[I��q����ca�1����
d�ߥX�|[�*I#�o�1	ً���d2�x޻Q;�~�p�VW���19��Ǡ~�0��ku�'����xQN
WD��V@�,�WN�w0���T���v,�|�R9Ԃ�\��]đ�Ș�"m6o�0>2� �Q�����O
*���iܷJʘD�S��D����oۧuq�L��&��zԃ��Q��SfZ�<���#&�����"�Cn=AB��N9����]��V�x�����K��g`�'�M)�ĝ�v��������[\���d��G��9vZ7[M6��9ҍ�Ƿ�VҦ�J��"&�MT�Qͣ�L|��E$<�����e�J�(m�T������ٟB�6�@�����eÇ	ܔk�K&��S4��q>h����zR�6H	��M�9�j�t�������?���@��YXg�b
T�(�pv�=n�v`��k�ǟ�Pg�S�e��{����/�o�9�:hA�O������i8�)�>��kK�/<t�7�EqMJ���6n,�2���!�ؙU�:S��u�&sA�oE���I��r�����U�č�^����Gn ��(+/{$ fۃ�a��f�<F����k������r�d���Q1���b:-s�%c������[d������Y�Y�L��[Q�Se�7\GI,�%S
:2���،L�;96�҆�@�$=�)���C�x����_"�X����ޭ[���N��&���%$c��#t��[ʬQ�F&��#�ckX�ʜ�_�fÞ�����
����=�cϻ���A3w?����1��.�.#�KO}����+E�d5�qZf:@: ����M�bj�7ڮ=�K^t�*"���1���y7򡉍��&���� ��3�(����P-r�;;�����R�@���AQ�����j׉�Ĳ�����%���+d������t�bkr���CT�l� BCx�\n���+�T:/�������C���"p��32�X�׺{V�۝��'5�	\���t���ɵl��r�ѯ��qΝ��,�S����O̶P,�Z�Z]�R�?�BJ�κ���B�U��� �FG�sJ�0$��7̯���-j�����6 �z�c�(��D-�U�MR(�{f��6�8���H�	#}i&��"e�V^��a�� (�^���,��C�R$�)s�O{��\���(�jT|=lg�Х�Zi���Χ�b@�%�ncnsLP�PVd���[4�&n4B8�p��"~f�Ue pXX�5p˄%�ܗ�N�h�a:��v<��D�d1[�9��0��6��I��ޟ��z���+C���r�h|&4��y���Љ�Y��r?,e���8T#��	��A���)�8��ō-���7a�y&(�kBFZ�]��~����̗`F���LA��֮���%����1�A_ZQe�x�w�9�y��p������99���D�NY��S8$�c�S�dp@ȵ$t�O�y�%cE�͉���ΌB���#_�q�����I���	+5?�qf�[�<���`ҟ�JC �5�_�v�y��%l�dD�u �޶���A�y�G��b�����r["��j���%r�l[O�J����-bg�Nrq�%ub�:4�ʞ���(��,�#�B^�pV\}:ZI/-tq���\螄��g\�F������U�(�vI��g��Tקghg�sK��J�J7F��O"D���v�>]��b(��4�S���cTtBqF��NY���⛳́٨�^c��̴
Cj�nU\P'/�/Aj�����0���)�N��f������d(8���l>YT�.h��5R���%��`ە(������&�`�����o.��9�^��T�9��*~�vD$ɽ�>�dw��X�I���(�r�:�82��t���=$/M�Y=E�=�2;�3���?/ˤ�`�S�Y�C�뇡Ί��.0Y�o����)7[tZ��|�ff�tlō�P����|~�v���7E�F�s�A�Z�[��~זĠ����8g���!
`4�u��]��*.�{�R�aZ��;�/���1�u��tlْ�u|%�����3��{�N=C�X�)W;�> �r\�����M�k�.@��#n����c+,*:�	�i�߭+����&�]�8�7
yo���<����(���$|Q;��Q�A9�,�͵1�1���Qav��JC`��>a��㺒ø	�����{����4c�\k��X)~��>� �v��,���V�A%������RX�*�,=�ꮩ/��7R��A>��t��� \WJ��z��R�>��#%�b�9��(�=�]Ёv�,n<��H�
	;5X��-��'��#�}�*2�o�������\^��wOC�ʃC�B.�(�'QX�`��2ۧ}����iR�B�u� Zd�R�fn��+%^�|X�%�G�\5�<%?��O1b	Әr >9$U[P����/-yΗ'�֞�Ү��fd o&���[������q�"��GdU�D������(-t��S.�I��/ㄭ��d�,�C�tK��gE�����#"	���19�`�xc�)��-�i�O�y������>6A�j&�䦏��'�bк �v���H<M���!����+�I揋9���q������D������9�~V���T��c�:Op\���A�S��9��-��~���^Wփ�F�L__~^&���2ǂ������9��JK�^�*}����SY6]/D�i��t�^B6��

�B�ݗ����](*��u[���Z�g��V��*���On��>̢\��T3�q�5���OcHr|0T��p_��+����O_!K�	�o$} )�9�*Q%9!܏�n�o	*�P�)=�I��H2�4�P��\�����#�ŕ�"][�Ť:E4���ޅ��s�̃|B����+�,�2PԔV|ߺC��"]���_��k�mО�ZTbP�NΤm��z����2��&�<45N�_�o9���3��Ei>X��nB.HƤEV��{
�/{r6
{鄗<$B�����:��f�q/��2��A4�D�}��:�p��I�Ҁg��JNE���Ìl�Ar��-[�)w�F���z�� �;U��`�i�$mW�j�)\�~��u3�E�7r1�8�R�o�`ڹ:Ro�~�?���Z�u��X�d�4Χ"���#�R�_W6m1I#���χ�R ��s��b~��lX����@8y�yS��j��7����z�:�0-�7m�U���8U��F��n� c���+�#��Cs��Pl9��k}�]u�}ݚm�N�s���fC�c)պ��\�;�`�w��-�i[Xo���3��	�=i�H?��i���վ
lñ�9��5ܰ<`����藭T����0`��_\h\�����=6<��FD�W���D��Ӓd!,�D��v�MnCO�PM+J`K��h��{�	�H�w'��y��%$խ*T6% ��"�X>�؁K��2�kJ��XS��iD���CR*,�jM��ׅ(����@|����F�hF���+��~��WJ��[_D�B���r�xp"����X��`p�������j58v����dߍn�(`.�G�/�����̂�=q�W���~C�*�0o ��:(��1�B�'cY�l��$�A�[��7��F��}C-�Ef�� <���7=��g6�do�_�}�Ͷ�z��;v��xj���J��*���=6 vҼ�F�݌�H�AR��FRD�C�l�(GH2q״�Ľ���`^&~I����3���ZA�NM/�,����0�����k1k���C�'L����㧁TY�v��έ����5�*�C��*R𰟢��O��Sʊ���N�ʐ�c���\!i����0 c�u�`m����v�0z�q�)��_��̐��D�V�Q�-�.
���|V�p�:� ���Ҍ�&[�Q�.˽dQ����}b֓�I��К��@�w��C�]���>>��>�A�Nxq,�d�Ӗ���@)`�$GP����S�	@�!^�)��*]��'���	�ݽ�)��s���b���TvFy&�ڐ�o����XqY��P�mz��l�<M9���g&���O��|� J�(��l�K�6�SE�|s&R ����O#D�ó�*����W'&��z҆�߬�K�L�As>���y���<���
6.�޿v�����~$���>]�Jz��0�g_�,ؐd��!k?*��`̌�	�@��,��!�Z��ۅ������_ܨ�mƚ��\)����w �7�.3�L[O���zks�=��cyo� �����˫�Wz1�x(L@4�ףMt 05��'p���o�/�{��CqR8�=� OT�c�W�j�:_tVJɌ65�M"*l���7�	s.s���A��=�g��Z�f��,�2s-g�W�m��dg.���#Å�Њ3�'0#5p14��E{��R��@�	h��7�<��� -J�H�q����߾.�4����c��ڜ� G>�k�ea�@�eH3V�Dk,a�b��/����:��s�/-6��μ�:Yf��-�dw)�>T�/_�y��^�C/��v�`��)����>���#cJ��(_ă�}<�� .W���z��c�����
N9Åט�ת�:� ��&�B44'���Yk+eڥ���f��n�-���$I�G�O��v�8�f<�ֹ�K������f���i�����ό�atB?�L��zs�B;ȿ�@��m���D�=�KHλ՚�-2���¥�E���`C�����u�G�.au��S���I�;|F�X��Q3`�nS�o��+5�:���A�q ��'�I�l��W	�E�]��,y�Yg,��{�yNα..sO�Z�C��/��P6�%ަ��9�������(6��aB{��c<���^%���0�ß��7�LQ��1,d���+�8� `��q�EN����V�� S�?@\|1��I`������񓙹�8 �%<Kd��U�j��.b�.�G�e�ϡ �
WsB�{|�c��t�:���Ơ5`�|�u^U��E�?�
�2 E���f��n�����}�g)J�������ۜ�á�xV�Ɲ���b0
H|bs����r�qg6����+[��S;� |;��&��s{?/O�ܣ��PC1{�g̽e���FK(�}?B����~�H�i}�^���m�)<�)�5�r�ÑXsy�-�sI�j���J``� ��H{2Ne��HxϾ)#k��&8,��r�>Y��˲&�މ��
+��~���ֶq[����X��`L2
=����	�eJ��s�(V@l7����9,�����8�߃�`JZ��a�y\�3Z*p>�il����h�2z' 5#��\C!�2�/���j�C��&�؜=��^�	��E��O���0���*]���r7?]쏞�`�mޖ��H�bR4��Q4e����m���;lg�!��������{�LF�E7Y_owL��Q��D��:�s�'���&a���	)-㸤�b�b.U�P�d�mhRz�܆N��(�2���٧V�v�r����^^��黇��ՁFF�@���X��$��~#Dt�|�^Ca�?���@}Vu�����R�>��|l���A���a�c'D��6�`�t��᯿���us-h�(��<��Gk��n������ۯ��,R�xc�k����wpI��`��f/�ڋ��I�(�U��;�N%�F�;��i��M0���Y� ��ߜ#QI� �{z9�0�
�GN�r�5��eS�J׷B9�zv��C�	�*�����"p��Ua��_�7�k%`��=8;ne��Уw5�ŝ���B��9����nݲ�̜�zx�Sу��T��g۹S��h��LC�[���A��|�!l  �bf��!T+Qy�巈ֻ������U�� eX����G�Ё<��˲X�XL��'D�m���}W��߇���i�� ����pm����3�U²\ٯ�X���R]T'l���E&�!X��Z�;�Bs��E�QY�۹�X�9ybM�����cI��lG�0P`�#��fB��!�l]�׃���j�(�`�s�)�g�/�4��~�G�p6�2�o�W俵K��ag�����G:�+<�Kӏ�E6�u	.�pˋ9��2j�]��gO1'�����T�E��a� !v���WÞ#��bqް��$�H�2,*Ko�������'U#Z#q��ivE;�"sս��tS�*�����Ď��`�, ��F�鋮fmBL���~Pi�(o��F��V%�p�a'�`]�fU��Z���A��@Q��K4�����\�e�m�s�Ѿ��~�wn���D����v1��#�%�#va��-_�{rɲ��X�d��Z�Z�;V2`�|�	�l@�(Z֍4#���Y<L?2ד��3��o���
���TOKc�ꏯx�E�L��P�����M�[�Ŷ#\�NuBcp��jg��d��	�cIN�;�)�:ߡs�{��)���vV��
H|H
$���y���o���W�m�ގD\_�:�chK��ʉ�ճJ�ŘR�5,���U����1��p�����/#j�z�3�j������ �Y���GHߎ,c@H�4>�^z)x�@z*BA�X!K&ptKA�H3ײm��i�w۩)"��
ij��6���1�m�]�?�H�+�@�z�6֜�0:��re�'��E��:�#V}�×#h�VHT*�#0/tV颊���Bk�ag׭	��Ν˪�FH���dł0އD�PS��lJ
��ti]������^~�mc�4�ऑ9�LF�fB�-�`���$~�.uTMi8�l�8k��xb�(�qh�4t�.rfV��a>��y���d>=�tF���n~b[(��s��#�����R�>��5�S�ܗx���N�>��ާ�o��$�s����]��nq�z�f�X^��2��2b����{�g3]�����w�~k:)�����S�q�'���US�L�ī�d~ɱ	�6���B,��A�!<�b�p����NV��VIe�*Gy�b!h�Xe��虛�k���`�pwa8��b��/b'0����8�E����w9
�M����G�p�m�Q~��D7%y���~:�;���,�S�9j���d@�J�_�ώ��y���%W�vIP����\�ȗ�]�'c�����i��.,M׳o�������m��X�Q�#M��ܣx���e�h���Sed'	�%Y���Z���ߜ,Zv)
�l���Mň?a}�ڹ�������;��
��"�X���ҙ� ��NwLH�Y����H�lE�aS�����hQP�b���&򹃲-7���[�����*&�?و�����P��0s4ᵃk6���������9���	���$�&��,̃����l��%�9���L��0�rӗ
�ĉߏ#�g*�lMH��ύ�W_NH lB���X��f�3��b���~;S�E᛹�"7���<�	�(�ֹm����&�����O����?3k��~l�b�"y.�����ד�ʮa�^������ +wSPC7/�;�N��Y(j�zy�(C��eة���R�����+�x����BfBbW4�_�C\���lS��lonʓ�-)��2�r��aTb��A�_s\ ���\+5���q�U5'���	��a�DA�w `=J��0��@�(Dꩊ�jM٤s(�V���N�A�7eʊ'Q��=�r�:�(@�N�c�?�x���?ñ^Y�ȕ�*Be&Z��j�QS<����Z���#r��b�޲9R���"�p霤�\��tS���-l�6с1p:�/�0�$۴%.�-�4�=�lz�8`Q��V��l���'�:ɫ\[�'���n;�U�t�7u=1X��_)ǭA�۫Y��Y9��mO��VNSg7�� �^Sdz��_66�Mw.e�B�Q5o�G�2��ʓTG���q ���Bg���%_��<XC6O[����f,��m�����rU�e����Uk`��5WW��)C��;ѽ�6��0��=}H�z���8��w������x� �ON�sRH���@��*��a�f)��0�$���9y6G� �	�������V.,�ɜ�:��}ȷ�A��3vOv��X5�@_k.d�Ls'�o�0,�I8����R7-��#Ę������j^cvp=}�di�2�n�ۢ��Nmm懠�+9�� {���:Jc��v
�vgPlRW�d�H�ќ<O�p�$7���ɛP�����;
��W(�z��l?���Uy�^Ց(=���̕6��p�y���'��E�D�A��B-˙,��_Nk	�RK�2TH�p��̕�U��Ҳ��������q͹m<�H�IM!��H��
4>WZ�1�K}��U�]U�%]�5�H?5l\߸��U�jB޷d_0I�=�� ��5H�F�l:$v�3e��u���Q:�:�W/���x��û�O����,�L���X�<��iw��d�V.T�O�.���ґ}vN��Q�m,�%A7a6! ֱ��!3��L�gsf��d9p��쬭�w�[�����K���do�]Kz^�]R���S +����;"��Nm���@o9��� ��{��ڟ����D�v�����c��i�$�D�:�	��T7u����t7c��X*��!�D��>��ҳ�DY�������,#���O	װ/����s�Ō��ɉ��.���Sz6���6�j�^p����8�ݏ_��i�^��1+���� ;cge�*�څ�y=̜%��$���K��|,~����Mo��~�?o���������Qa%Z�P�{=��GR8D[?�z]r�^��Ejż�feA&�}���fiA8���8����	Z<���(m�E���pB����q/�z�V~[�KV}?����	a�m�F���i�K���W2�_A�2���4w[�p%!Y�Mֈ)6�	H� �ߍ~�?��9s��� 3G1V�����J���Kɼ�+�Ҥ!��b:z�6��V�t�r���^�OK!��6	'^�o4Y��ޜ�r	��X��͢���gE|�����p�*�j�K���`IC�B�o�?�X��J�2J���v���G�f6����uc����/��M3m��T):�e9s��"���W�E��3��7gI$����? �'YݫW(�A��W���Gg�����8ҭYo��R�IReQb�qc� lXQ���wA�;G���߾#�X�NZF���i���Ĩ�l����!�*B���5@?r�R�y+BJ(v7]هF^$X;o��#m/����M�Zy�4Sb�a]�H3��Р��Zy�F}v��ln0�����;�t�8_;��ӛ\-8a'���/��C&��s��NW�B"�D^��[��ܯmg�Ny�4��3H���>YS�j��Mʑ{�\�!���=�������_z!t�1"`-�4&��x9��&����j'�'{��j�0.Y[X�0O��P/�gMy�^��-Ca&�Cj�b�O�����R�#��,�6���Q�����I�9
�J�z��d���{�0*.�\d��#�����̰��k�H��G~9��iP�ݘ%�'VZ&O_�0�y���!�y��'O�f��(T?v;V[>�Vh�͋��*����̕����u���	��p9&�"s�K��c�ΠINѪ>��F���O�����+��O!�y�(b�L3�\ӎhL��BzR�8�,����'��>t)_ub�����|H�a�p���TJ����ܟb8�V�PN5Qy�
hc��o����H-�F�qC"�~�`\�LO(��r.�Z��$Ƕ��������335S���m�j�Q!}������%�̴>�-'�Kf?hEC��i@�i�n`%9&����ΉT��/�n{�bI�� �s����rd�|�� ���0���Ht%t�&��=	>8K]KJ�g���TK���fvx�ŗ$�ڛJX�%�@��R��#�����G`
�Xzc�ڗu�x��X)tUM�P i`kf��������JT�@�¡��Ϭ�΍�
���1�,�<��5��z�
ۗ�y�) `���b|�E�?�&��2vjV���+(����U�@��F�ޣ�,��ܭH����fR\
?K�$2��^:bV;h8�Ǚ���qP��y&f碰O��]l���;��(��t�U���\B!�E������%	� ��g���K�*Ͳʏ�E MqK�
�AGH�v_�g�N˞���!⺃o%�$aB8��R�������6��@biA���d��۬�2ʍ����O���%��ub+��E�q�@|NG�`�t���*��RB���zS�|��Ş$k��<)b��H�y_OZ��ݓ���^��v�c��0#������%bz�1��n�1C�,��Ɲ<��H�3���;0��v����,���ь����H�6?�j�.� g�A�Pȉ�@�_YU����nvGe��w5���c:8%��9�5	���xx�v�5Q��c���}��E�
N�_�|Y�*z/W�]�Ʀh+2R�2"%wyyS¨�p���=��,J+:���w�`��L[Vd���%����,ɼ-�I��M=0�� �c���ۭ:��s�zH�$L_�8�L���	(�i�]�ʫ^��p��9D�yq\�ǒ��B�_R|>K�G�'P�YL�V�Xr[t^�S�Mb;��=�U�FՊuCd���]�Hb!�ilw���Pk�K���|D�4}E�p�(n�d���Y�o�)��Y:~�fz᪻A}*�jv�jؗ��bS
=p�_ۓ��~ ����'w�%��GC�w�m�oeF��AY�`������� sZ��l�����\-�j��LG����n9��)`%���1e.v��ӭ.�-5C�����B����@k!�"�.1��n�kK���$d.�P�6$�ciP�G�RG���%
��2FRk.h��e����J|WC�[>ho&����`WG�|���6e�|�#-�jnwW��I�+�$���o%l���j�W�Aw�Xxg����͕�-�9�z�~�j_�_
Rs��){�ׯ)T��*ՅG|,w�������kd6ٜ�*�`�c���,���[����)�H�w1c6�����n�����2��f��G��>s��|��[O�dʶ�Z����Y\|����Ҏ,(z�HbR J��G��u��gݐŠq2b����B6�Y2Z�5�7ΜҚ�5��+� ���j�u� ΎzT�P��[;���v�L��Cd<��5%�*�N	SY�=�U�-��]�i��"d�:i�v�h��	��'TOg,!U���Vҫ��Y*_���J`%��B�;���c\�K+)%�7�q��t��_�ORs���^�7��{:q�v�QڂB��3��������S&%y�o��y������Y=��s��g�V�SX�g�0^8'bR,-�Ͼ�����B�w?�\T u���?��ZƗq�Ġ�s�b�l�]{`i̯�{����gx�L��.#��"Fip���l� ��v-j~���ڦ������>?�NAe�O�J���D���.YK��ss�
f�Zt�8�Ҏ-�hH	����׸�e�m�D���T%���1T}�$d��e�߰Ћ���;t�S�	g�8����#0��9Gd��X��d��\ж x��zy3����L'�pr�)N�.z͵r�vx__��a������t�;)�B�w�_�.n��v!ı�@Sw
�f�N���dKX�Q3NB����<q��F��Q�U���sH?d�7I8;��1�*�ŔD�&�TԎr��W���y��6��N{�sj�R�`I"�K���5�������@���<�qS����8����0�S~����4�=_�I����e�;����9>�0+�i�]��R�F}x���A�ޗ���s�3r���� ]c�i����[���oNj!N� ��*�����d��jEG�b"�}�$7�:-��=��Kbq��'t6�g����rE�s�,�$���3�pR6��*B|92-��Nt�FC_ #��J��
��Cq�(g��-���C���X�|���#R������;��ZH�G$v%Z?[���j�5[��� �>
$^N_&my:A�-������V���$���������\Ov&[.7{��L�"*����	�
��.�Rаy9�s�&cs��!����ۻ���(��W�{�.�y4}Yk�K��lbh��܆�F�7;�'_!tM�˶��ma��'s�%s7��#�d�a�D��7Cp��'!C_�(HH�&��tك)��p�$�L�C�f��o%�J�/����^� 2��T��L�w#�"0ۊŋ�f���aE+�[�N�1�Z��w�
*�g�1O�L�Y�����fIʣ�"d,�>��z4K�q���k��=c"�� ��+��/49�Æme0��:qe�ג3���	���3�d�<�D�C����Y�:	x#��X�\nT6f٤b����]�S�<�f���C٭��ԉ	` G`W��)Uc=q�1;���R�O�
�%,�ј)�\��o'���2R��*�!��]q�쯥9>�FL��l,�Vk��t[Ԗ%�춾�I
�_�.B\P���O���ƃ"�0�@z��+��6;���c��+���jµI$3�aDAO���~��k��B�*�j�)vtYb����9�`S�y�#F���6�7�f	��($�^Q�+��b��'�~�ϫQ�l+|+$��JPݭe0��*6����F�x	��z|O�'��a�����s1��t����]e���'��se�n}���ܾ*P~Y�_�/ >�/?.�����\C@m�1���߅뺮9�z�����ރ�r�C!�<�AW�����,�r���z�N3ד�AXi�,�΁�.M�'��w�Қ�wm�4�
Q�m� 	�HT�J|ޠ��n�Y�����wC*��/$RlD!Nd�c�~������8����]�E{m�jf�8�)�Q_�}����=]��.��mJ�3"�D�
Ge��R����a�D p����t��޶(� �t�`I�����E�q��l0�;��������A���a[��$��*�_f亿n�]n1Кy��F�:`5��&�|�^X"T�esQj���<�?�};!!���D��y��ט���x2�Af�����2���p�ѓ�$@L�	R�{o5�1���K
���xy��C�t�{�4�4������x�dm�����@�S�P��@=�LF�*���U4Bǀ'2����d;k;�x���2�Ƌ� ;qY�NB^��pD����Z�����?:���8��Z���{�K�,B����c��L���������E<�Q�9��·�UQ���p��7L�T4"�nU�!.NE ���^����}"���zI�!��K�����T�y؟][����|�oC�^`���3k�Yg���T���c9!Z`����
��T8c�L]\��?�����!A=���L�g���Ρ���~�Tj����;�,W�'Z��f��#��㠍���x��/��u`����P;�̈́<��"���?���z|-p5�����;�r!�d�~%S.G�Y�� ���)���0j��$ɗ�lx}��Q��ծT�F����[`�?�s����r��w��[�!��k�D��R� �������n���ڗDq�2R��}��gd��p�m��9�E���B�T�ȳ�ԃ^A��7�1;��y9�����/}�k�pGȰEθj#3��h�P��@Ǚ/�����|����G���;"X�=�v�kX���<����G$M����%2�m�d��]�`:���'�Nں
� �Z�*���_A?��߃ ��kn��V�I�#��b��꿙o3��1�r���0����#w�mX8ÎV|�Ir-�Ӄn�ѡ�ƚP<a��5{ �hAD�|YK�Zȁ�i.V<o5f�6f����y�X�}0�~����q��`��_�0��3:D?�t�w����g|ԍC:yb��~����}]�_\�@�W��L�j'`,�pu��I��)�jp�M�8F�|L��n\������gu����Hh9݆�߅8�\��l1X6|Wv�����`ㇲ��[;�[�P�OQ��҈���<�
`}�$�@�^�f�_��͚�Łfn"�zj��^�<���1;7��c�p�wʬj���½}'�R�u�tB���ا����~�,�OQ�*>l���I{��M���ֈ[�v�t��w�����dׇ���m`>�<�3;#���̬ˌT����=J�}Ѩ�.��o�h.3��n69�U�b���K佧�8�jt��9�q�B��EqY�P�/�h���_gZa��wZ�BeN���ܰ����Fb�'C���i���<</K�W�Mī�"Սi\�XK�>��Zv�0���;c�!�!��XI����(�Q�y��Amk��;�:_�1��w����a�������Go�{gB�35�\��Cu�����&p\�f1rUN ��ꖑ&i�.f��f��ٝly��.w�m`��@4!�jy-�bi��R0/�nO �:ҭUr��ORIu��י�0�,x��0ǵ�Z�=k|�f���턈[%.eW�
�
�;�^yV���^&�v>8���e�\�hc%��uF�z��{������5�z����egz��Ϝ|��U��jm9_nx�D��(�[��eN������� ~�c�e�ķ��j�ZI[���iI��8D�#�a�)��wN�h�����\m�z�^൲�Y���,TP	������7��a�������KF<;��Ū���<n��q�Ra���Q+n�[!7^	 �|��}�F� �b�6��J�l��i.��#�/�#>	@��C(P�R	�����YlPġ���8�֗ܝ�' �]����[I�L�uՃ���t��9�{%�l��j��J�H��V/uh�`�ڟ��h��]�(~@�7�.(��,/�{Anm�����^�f%��N!��#�%n��@�M�=����i7��X2뉒Md�Sb*���()�ԛ��1(��}���T�Q��#��b�J��_�Y!Uu�GXv���e�?�� �@t�n�I��s�Ҡ+L�M�����窽�����m��7��1=/���Pl���3Awr'�ƎUDB���{�y�_�x%��Ȋ3#���-�tz�7�l�}r~��j�%� �ѭ`��¸^�Jf��ӨKs��̸����#���`^�D	{I��m2Z����E���z��)�����;��q�:e�t��ufs� ��$������ڪZ#��cj)6|����\��F��Je�RQ����Xr�K#��J���/o`I#;�`��+k�d�_`P�M����!�^�Ig�\,f�/�A��)'琗�CËD���/ye��Cܥ>��$t��p�p��+1Ek҉�5��@��;;X����d�C�m{pi��������"ᓙ�����`�g�|^����NҫҸ�RmU��CF6ՑIF�,���]	ψ��\}L0�������O��&+ۤ��o�ۊP�e|qx�v0�8/�j[0AHD�+�:�����0HQ6qv��0B��J��`��E~��rem"�ᄃGM]��w댼�ɱ�e	�]_�$��#���d����┐sqn�֗���[��|?9t�򷠽H�]����m_��O�sW�K$10 ������s`<�����wV皻�c���z4/Q9�f9�$��[��*���j�[_�.mp��kz͊7��M�s6�Yj:SVɈ*��'g�U�!�ޛKO��^B���:=�p���Q.D y�=�(����I�-u�a�~��
Rt,67��������S�@�B?�#�O�_��y����S�����4���K��/��`x�$�p��`��r���y�S(���)L$J_�,GD�A���R�O��a'�as_�pbS*�ُ�����3rIs�5$�5oz�;{ I3�� �e��>��R�o�nL�5�Ő�r4da�I���x�����h�_���c��ϟ�d��ɜr����Y)��bѕ�9'�Z�"�ƨ�d~������MHݱ� �(�#d�^�Am���J"K.{|��"�����tj7���(N�BT�r�����a�~S���*�<]'��s�Jk�H��E��V�ۣr���sJ�4
v��
H�Z���%W�>30�i���X>�Y�S��%0��m�%��H��賾���l���u
EQ�͜��{ W�D��-9�����d?|vg7ք�>�|w(�4F�n�ȑz'��u�1<�,��E�0�(6.��q�ҹ�5�i�O�{���,�Y���{G�\�����՞���
��:/p��bG�	�%�bA�{FC���嗟�Q�q��ݲ+�F,:`���5Q�0���y?�SN�z�~���3�C���m�E۔lۘf.m\��i\d���8�r��"��j����z�G6U0x���8��8��_k��0R%A��>��~sy����OК��<�uF�6�ؔ�x5Y+1q#@�Ȃ��3��Ƒy� _���S�_����x�r��g��ƿ�c�E�� ��NX\2��'��jq��x��N,L�'�A��X0�^��{�$�c	D�zͰ��B=6��[��&�,[)C��T�,��(�ryꉚy�x��*6���Ͱ�-��1^�)W�v��m]4�Tb�a��_���G2�/�τ	��H9?����kuشKN�Q���$���E��塇����1�.N�L�t)+�g��f�&�YD�|�i�� g�Cʉ���A����z5�e�Bu]l��_&�,௚�*|	y�
�d ���̏I�6��
��׺�=d���#}>�b�mؒ���!�f_�N�G�1�������|`�R�,3R&c��9�ݯ$�c����i��C����C4��L�Y�N��s��$X �h]�O���Z]���[^���K�K�'��A�y�#��y�8u��tZi�C�Gz{���6��;�[Pq�C��r0�r�m����[�ѩxIcH�Ӽ�6�?���K�VJC|s��:��u~33ı�v�4VXna�Em�;M�����Lg��ul�rq�aV���v~7�7
��x�$�4ָm�����K�z&>�Y�x�:�,�����Q#�����储`�$ G`�1�@�r1#hܝ��r�0��c�H_R���yI���.��E[T�\��*���r�ތ��uZ�T��X�t+��~񸀎L���te\/�7�G7t�"��/�@JB��$� +�P�_:�w�Pz�w]�K�f5Siǭ��.�a"Do����y0��D�A� "|֭��Z�Y�{�����W6Ο.v��7H��h��[B�r��*�(K���{������m��KB�<�(������g�p���/>Vg�#BE����йPקWC#G��6������0f����)X����Nd �f�v��$2]'V�8�S��`�׳f|6������N�hj���+��1?T�؍XZ'���p��vf�g>ϊ�f��]�k"3n���K����u�f���m��?uCH7��.OV`
��	������&ޤ%E(�|�k�1pu��s)-�L��ro�}A�7q�YzlKd�0��Rz�A�l�n.�dM������?P�T�Q�;v��@��D��KqGh���~��`�s��͡J�8_�E������������m��a�=7�(�:��Z�T �M1�kӟ]���pjޔ|j���X���c~����R�$�CB��O���|s%������}���0���f�%ޱ\~s�eud���<�g�*�f����9�+0&�R�W��7Յ�Le�L�/���7y�5`��WF�*
�.���&V�U����G���v��n�!-�BVb�Z,:d�ف��.�D_�~���W��޿+�J0�|������� ��i��9�Uk/{H�q���&,��sjC"Y�U-W���G`B-��1Ż.Ј��SQf��(//	[��b�.QY�|�q��!��. a`������y�6���M���ʡ��}`���?=�I���i=����\��-M�k1��a��GcA��R�%�ޑ&�=���?���U*e��?�o*�xOP]�mm��'��P�g�U�N�{Lʩ��s�M�^����Y("���X�ʵ�!lV�ي^����m/X#���P?�n��{�����2�" �qtjf��G`0?�.}������1�e�e;�Z�QUJ�!fs�}���>��$e����V�q�b=$��;���;���1��{��Q�1s��!q���)d�
�]K��}��Z#L!z:DW�&*V]����x[ظr炓�f��62��
6�ӯ��T-�k�`D�}m�&gC� ����G��@���Xad��e�29���.���M#��SȎ�AԦ�C��b�E��Ra�0�T��o%�lx1?V���W���Y�^ǽ^΁~��*A^JH��Qc�����ѵ���1���(&��Ν-tH<��ճ�����WY��ߢ�@���n��4ͨ�JF�
�p���׬����Z��b��2�un�x��g��b9[E���F���j�^��g��P'�#�5/�1�A�.�G*3��T�d�Óy�C�X�ު�`�<��/fk ?����?�m�i9�sx�R�2Dt�cyq��!aك`�D�uR���*x�bZ��İ%�4����D�i=�'��.�z=�\"ټ3!���	�̏�m���P������V(Um�7V�c��.�$�2!'��S���d�58�:u[��ŗ7Xn`�@�����2��봋��K�.շk�� /L���:0x�������K8n)���.�)W�^c�:xO����4�D��+���Wȣ��Z1�P���z^(oQݺ;�qy�m�Y���/R:oj��Ԉ��8������%.�ivc�ߏ;�{C��8�@��]�	"�K'�r��b,{!e".-0��)>����m����]����%!
��ӟ�����9��[�D2H�:;WD�FWP��u�3��M����r?���D���x�z�E��Å���K#|�c�L��V�X��=0�����s{6+�2��$��VԘ���'�rv(9+�=zh�k4}�D��=�K���ە�:LA�8��c�#j��&<����GEW�u�(J���O����\�6!-P�Q�`�t��ߟ������TrZKqK80�8V��~G��DQ��(����^w��U�qvNW�G>u	����.B�ën��RG���n꿶N������VL{�`Bv
�ݜ��|��u� ~7�+YT�{�]i�
r���6���h<�O���ERQ��(�}g,�+9�J�����\��k�P�W� jؙq�e�?h�L^À�o���N�6P�jG�vi����2fz ��~�6�2��	����[Ɏ�סg�"��,	g�|$m�֓2M5N������\�P�"�;5fR�޵��f�T	؏(��0�:�*��K��'ψ�c�_ٛ�Z}R�����GɈ���P�ݨxi�M���ߓD|*?ŀ�L5�ƒX�s/���k�	�Q�)Q�F��Qϲ{<R��*#a�OkL,�]�mN��$'I",��Gg^b�}���+��Չ�S���RJ�n[�5��@�~�γ���γ�R����d#�R�p���1����ݨidM�z���|�Y4M����{��-bL�$�9����|��%w5�~��q�g�^,=�i��#�m'Om�g[.��kOWg��h��>��O�E;�3NvB	L��6W����ј䷇��K8�ٓ� pd�����Gב�ru_Yp�ь�"�\��b[P����DR
��PqG�jo��%W�k3&׿�c��bP�c_�g���!E��ښr�#�Y�صü����'�l3ؽ�\IK�A^,�
����(�"�p/�!���?�y�������#�9.��&����<1l)\�����%�P��6h����:3�^>�Z� ]܎�=�P]8��Ƭw|C������h8�T��֯�4l9��<#^��g�U�Gy������:Ln7�i���{gE��懪�-� Y�=�'/��b�*pW�}�=`v������f���������ձ��B���R߫d,d��<��z�	�^vA5bhT@��k]+7�`I�Io[��T���vr[��R*����.�	������8�?�k٪�����	�^B�l�SG�����>���c��U�K��>Ӱ[eJi�O\��p�15�s�E���@�GO{��	b�a�Z9Q�b�L&b��)��2$�K����(�ckd�𦔗و�.����wݸؖ�TcNO�pG�*>;zؔx��2D>�������{�딜��h�����9}cn�6�J��ߢ
8��A�v��F�\�<ϸfb�Zne�(?�F�=%&Ũ�+#ሤ]3c�8�{��i��t�j���dn)��8?z�ƨ���QlxN^�P���]�V\N��X�dʨt�a@:i.Y(��Q�ۅ�S��Y�֯�H���G�`���}wW׊0i��x�Gx�ʚ��]���F�	�hs��2��ͳTjk?�Fۻ;\�����A!T��`����}-� |+�q�%�2�ѽy����Ҹ	�d����s�FZ�A�iQ$�ŝ�B�t��+�>���-�ߋ)�Lm�ᬻ[�l�c�Z�`:~6������߃�	��r�t~�۝��܁�'�_9nՆ.�?��x��0���3�>{7�o��"∉��t*yE�ť)A����SB�'n�c���Kqݽ[�AMf�}��G��p�'r�\.ݨ�#��3爃Yzhl��1�|��FeT��Gyp4�<�J��ސw n
��X�q���ڹ'Y�a�G�T����֯�:�ڀ�KEC������7�1�(nhW+�yY�q���;'_vXql�+D��$ �.�ϫ�G5���0\?����t9\a��N��yc�+s�^�����\E��>��/�G�HՆ��$��IX�~_�R6���=�M��a"�(�8�����i�7R l�@,�e`�!�=��ҵ	�5�U�g�
Ec��B���g�}!h��N5K�*�l��P�ӏ�)5K��D^?0!y�f�#s>�Z�'b���I�ZC,�m,�������e����-��*��P$g�]���Q�+����x�~r �.Zx��Y�Rn$��0iN���C��@nGG�s�S���{�ؓ/��RP�s����󸌵f�)a;��?ٞf�1>�,O4{t�L���?�r/4p9����ur�(�MKXѶ��8��|�L��g/Nt���+�o�qM1K�O�^�G	ثPn���� ���O���U������?�'���d���YŸ����M2Y4�d����v�kf�6��M��/0Ý\�N�C$���k,^�?&/���`�,��-C��L.�;S%��!�����5�wCO����1�~�/���*]�;o�*�h���%V�0�u�g���S�L��H�:"�2!�i$i��J����uK+�X����K���oj��t��}�<XR:dM#�ݣ$�#�RM�4n^�OC8/�l��x#�|"L<�{��-���A�ﺠ_�=��yщԏ���BM�<;�?�:���ʀ�5����q���/	��=!Z��`�5=���B�V���tK�8K[�xi��xS��4U�$Mw�Ѽ6\u;��m]ڕ'.U��>��H����O�]�� �/%�pKz9Í;Ar�o�H镈�@��nɁ�[������q��9阖��?�oo¾k$����|��0��\���U�rb��i<���ˌ���]/X���»�5MOc���TI� �@�āɕS�TJ�PL~Ѿ�j�ǉ���STN)��L@��`�?�At�"��s���~��[��$g�K
����		Ց�Z��WX���UXNȘ1��I _���rs��(5�c�?\/dsf`�٥� �9|m1Y�V)1���D ��@���>�;%����~ҧ�K�%Us`��@��[U����؜�	۷�����UJ������!��UN�QhH�����lK
�rF~A���s{���������^���{2��+H����=󐍪N�$��obR�ٛw�r�0Eał���i�y��+��s��?�@ݿj�b.��3�L���d�sd�-�<���Arܣ@Nݬ���9S-�ӳ��G�=�.�W�2����[vl���
S�������.�l<����5�},��hw]S~"gVS�򛖌����}L�%�[z�9����9��3]����߿�/eB��zz��Kwv����K��GpȤ��b���X���A��̋�\3η���mJ��nˮ�#�[�T�L��|��%��l>�Wo<����8���(d��5��^ѱ��+�q	�&BI���1>�}C�)�}��O(���0���F� (ʮ=A�Z�ˊ-����T�D���"Vw�,+����ӿ��������kNT��k�\P�� d���I[w�i�Z`T�x�� ��o-���	����|�����c�f�a3]�L�Ӕ�e��?����%���/N�><�V�� H�9��`��8rm��)vTH[������i�w�0��0���'��3��?JBA�k�Y��t��2��o}��&�%��i�;8��+��5}J@s��@��,���S��3�u)z�}�����{�(�BI���*"���s�b���C��]�:�-�]phI�����@Y�:�T��ͼG���y������j	�HL�J̂��>Q6��-��#��7DEJ��.��+I�7_"����Œ�7X�Ϝ��e��N�}8;��X�  gC��8c<��2��[��.�ز�!&MX�6�Ch�.��뮓Cd�D��z���SE��$�q��R��7����%�������2]���D\~o��kG�����~��S�6���g��`���f!괬"�R�v���R���v}�¢j��ǳ&&�ApS��⯔�nϰ����ƿ���$�Ü��IP�{aLf' A���k ;�|�S�����)_A̔�F��@ ��Ok�76�nf{��	�6���,�5[��{��z#Wn�������/� �DS�]i�� ��Ec�)��pO%��k���x%��3kIq���&�%��H����K���\�yb�xF��*�mC��B�,���cP��3a6q1AF��^�"��2���]'-�_ZD�e@`��E<;�S�Xҷ���oov�#X�>�X������<��/:s����b�d+���
v�֦�u}�|˸guΐ��X��ɀ9�򙨿/}BBN�'�ڸܟ�R��*	\5Ĵ1V�,9��3�3Zdz��`�֩�7e$�"�Ew�q���GQ gC#@�a<�Y�^�942 ��P�;��C�
s��\4rܷ�m��O6�	~':� ��&-O3�J4)J
S�Zn �s"˵���ڥtO�pAҔ��R6�4܅`�d��؄/�+)Ͽ��6U��u�������x�^�#�Q��xM�3����j�wO"�l�U��w�?��wZ����gH�3�N���hv�kDEќck͏)�H^���\�f��� ��Z��$S�"ҊXҕz>����o!����C�F��e�&�N�!��@� Z��RM��[���\�~�j��x:|��e:����Np��D�̆4�g��qE���=#4a�&�[��)0��c�V͖�9��t��F��L�}K+�"��IJ���w[�׆����)�0S+��i�13��'�����&��Ƈ��՞�c&�H� Wi��I�0��u�_V N�HR�ۍT���9<xʍCV�qf\�N���j� ��q�� ����HZ.8��Þ�$��3���Q����@��`�ʯ�Cp�&y�	���+�w"��eEAG1H�M��g%���s�G
d�R�ôS��Q9��V�Iw������6��]ظ���ev�)��#s�be�x�w�^�������LE�(����X�;����`]�v`�^�A���Iq��>d` �B�U���D*D��u8A�8�����L|���8�����9g�`�օG-����Ä�[e�`��l��ǰ-����I/ v�@z��;ç~��)�҃��&�`���Udc��0;��̛��Z�Ƃ"��	���l�n�`���d1&�ߗ}f��B�Ƣ��;I�ܞ�.�2x$�HxO|(�I��'=~�撢��b�"yh��	��$�m����G���ּ�6��\a�C���ঝ�O����+�_����{뀿)�>�À&���T�F��H�?}��|���墟r�gn�6�6���~ߦ)��8(�Q��k�<<�|�x-5�Y���N�h-�8Sҷ�u�E�KX�NN������g/��nF��c�+8�箛p'��Np6lP��#8d �%
p[~J^�P��>F��b��s �P��Gs��W��i���%��P>�Zn�}��W��QTSp'>��?�3����C��@��Ob�7ݱ�'��h�>��hT�}E�|�������<�A�3���o�T�68�����t!�WSaO��q��лL[���  )�S2����^�+�M:I���z�Y.�z�EN��"�^��z���K��@�Q�����ia-��)q<?��Bj6�LZ:�ڂ��g����1���Z"��-=7F�ގ� BW�[Q��(X�+w�=�!��'���PR����
�Iy��k~��>���aϫ�eЅ�!�n!
/ɳ�e����d��)�o�V��A_�C�RS��ׁw�,�%r�M&�̏�>���&'��f܊�4.������[Q����OpK�o�'iv�e�N.K��\��ߐ\m8;|�r�bÓ�9$��
i��dǮ���.��I��o��(Fc�UI`F1\&&!pİu��tH>����p�
>����f	�0]���J���P0�o�g���1��?ߍa"!-��VB]k�	����b#�"����e�N� Լ~	r�p5t��.�H2j0]�}�E��Jr�3�o�V��	�oV���b.؏4.��C1���~�R?�1vޥ`2�-h�5z��oj��ҷ[���fH�� �R�uv�5&ƕ��4�=v������`��Z�0�s�����~+{�6�{�v��j��j�*#9��J-�jЗ��^�M���3I��g�� �9Cv���B|��ZF{��HW�"���܊���UE� ���M�
*s��F����Q�ڮ3�rH�E��#r�������=Б��ߕIC>�w�Y�E��˖�S	������ ��P��G�!���D6ҽ�s|��Ոژ����?�cV�yfC�Օ�����Y���G?D3�Z7�qY!�
�� O�$Ȍ�wJ{Zt۹�Nq��&C��Ö�a mRa�P$�Y�,�|ݾ��T��X��w�<nw���hHU�(�#���j�\�Ӳ!�=gdНma.g#S@�"�`����;5�C��I�n��f~�9��C�ݎ������E� ��ܒ9����j�]�P2}�l��A�M�(�Kޅ�Z��b9����fj�C��g��Z&� ����o�`e�����Mq�v�_
��ex��դt�6��������<!�����+��Qw��bX����eO�n��)�����v+6b���&�C&����J�x(��0��p���3vl�1`�w��/��QP �]�*��	��q��j�\D2�Nd�L4
D����	<�	��j�ׂ�b嵎rF��Y"|�%g���N&�1�Cʐ�%K�])�H��H/ʺ�Ͻ�K�L���! /���=�
�J����?Ѭ<2$�6�����B��J໶LF��to6Iy9������E�Cl&?��]%xjV5)��ʍ0R���C���޻��*>x_�n��e���^:ְ
�&\�&a�|"r"k[s���5��m%�M>WX�5��Q~�y�8��'w�4�ͨ6ȂA��E��dT����t���*���K)�&�S-duz��6Q�}�F��;vO�-'ձS�;�q��}�h����L������IMt{��������n�O*c)CL�t!��Sx Mxx6!�(���ht��A�ٝ��KS]wE�S�b�|>Qי�o�c��DC��G�:��'^����l���7
�th.�����ǡ��^
��R'ȵ�|�%��r38���:\��Z⌙�J����J�hG�������tWuL<"m�3�!ܚB�<pz���T׸�Qz2ҫ���E+sF~�.fm��a�iaP�n��	��z+�}�j��39)/�p��5���re����n�wQyl`�
���r ����
[F������S ��gL{�̴cm'���Cu�P�����.E����"��h���KL�g:��"�y��vN��o�4��8�Яĳt��;A�����C���E�Gd`K��S��9\���X��q���gM{������� ��^�X���.H�5��'�㯚�&�J�����IJ�[��[���n-��g�5�b����c6��� ���ː�[�zL=)��#�cO��_��pBÄt�`��K]�2��np�=}�)QT)+�K4��X�AT�{P�0Z#~�r�Te8�-#a`��3���@�&���6�
!�tM4�z
:t�[�5:�%���/JJ.����໬Ys0FQ�.�Ă�SV��@qEz��
q|��n��ϝ����k0׵E�E\��%��x��p���P���Jã��J��[|��i���۳4�T�g����0f�'�A�|�kIV�tn�����b�OSZ���n�E�쳡W������,�]X�hֽ��{�H�����)�.%A[�PPO�Tf�xe ��(�\I݁k�d�UqN��=��i�.up9�W���e��d]{�R�����k�x�R������F�V�I5�D�=���Ͽ��IY�� "d��%���o��ɒ��qr�d.�W�>I���OTu_��\8�	g���d늴l���=�k�k�Į����@C�B�i�]ʐ`eL�bCg{�W�/���[�v�;�|p�?Y���*OQ>�{y�T��"5?\���b���.R$�s�����6#Q�!c͛���CLh�A����V��7�1���nk�����q+W��A[X�g��Ԗ��j�ܢ��kW�mM'!�f$�8�B������i[������C�1�f�+��xJ)�#��Z��ݥ	9S+��t,s"�}tǥ��E��/<�d]�jJ�RS�Y���%�Jl��Ō���c���L1��������R|�xK	�h,�Hw���iK��K��<`�)Bd�zx#�Zo,]��U9�?���p�+/Tl9���f$�\��g�΂���\��v�����"�R��̄*铳{�Qe��5i��WV�<�� |sޔ�4ū��3\�׃
W(&C��L�]�Ɨ�f ��Q���"z?����S�L:���QrЯ�S��k,6P��*���R1~��X��5�4�pSQ�y��3�*��=S�ATe�`.�ߌ��[�qb���w�����a�x;���j(��M*��W���X~J}LC	AN�aB3Ha�ELd�(Dy֤-�����dۖ�_$���o &t����L'����([ (�PhT��a#�v/�9��lXt��S�7�įd�3�|�����D @q�ԟ)_�`�Ge����*�����[��bjT��2F��sLr�kSp?�������E�(	l��i�&?��?~[�h�G �>93O����2��y�"ߧ�6�%*L=�	ď\"��A+�'���\�n�L�a�����vK3wҍ��}��nqeR\�xB#��i�X���z�D2�2D�ýY��Ax�Qu#�I��-�>�&�{�]l�����:s��F�d��qe��Y
����Lw�گ�yH���e7D�@������d��t-6�i3E�Z�3'7Ab��M^Ȇ�Ƒ�%T+�T�ng+)گ���z�Vf!2$IY�w���/>E{1��-\��Q�&�-�E�X���	;Zm! �~M��10�,!��P��o��
���|�v]��d�f\๝]��T^�z�S%Ɖ-����`�TnW�ƞ3��вZ�$t�]�L液�!��b�;�,�Z��
�Tܼ���r�������������],ʪ�-_�=�R��k��� �n��妮��c�����OK�SY�S�Z4�"��~�5|wM^X�Z�L;�ٻy���F���|���	���i~�.`�����"��B��E��\+��Yf�r�[<�0���6�]=b��.3f'ĝ��5�l�M���?�������~��
��g?�rJ9���0��լ�,?������ϲV�ij�t41�D�A�_�-���ld�^�[*MePpg�QO0Xv�B��o����)@D�]���M: ҶltnC�Y� �♐��lGE|�:���,��ν�>RA��c��l�U/s�cl�3v�MM�m�y�q�����k�w<��]�^�l�0��S���B3<V�}'�Ʈ��_m�!x(;g��!m�Rn�f��h4f�XA�� e����C����0QV����腦ӆ�y���Ja zƟ0�y���Y��)�a�50��Y|K�jh��z�F:�>��!9^P�#]�q���>���lRh�#ܬ�K_�5�ǭ�4̍���'Ekk��|�������{K`�C�Ao0�)2�ua�X�+0oo�|�#&�<�z�	�K/;|�P�I���������,��6��l-�`�._�T�Cd�%��9��Y�vG���`�U�͛�;ƲA�
�c��%�l5z^�tn����0��wc�ˆ�ǥ)����w��q��I��gh3J�����D14\���_�pC�&N��բ%J���2+cIR��*��+�:��֥|��[ݐ�c=��bb�F@���u$�� %�UE��9	<΁Iƨ���z�)2��&�t	����ȟO�).G8�/N�Z���4�r�S+ZI�0�N�
q0��C�����#Z����0�m�����J� u�(���l� 
��bzOL���A����9_�p<X��J�B2��-��c�d�(%uL�c��f����òS5����S�K��E�;�34v���E��~0��\��T�#.�k�á/#nV00����_ǰ�ZY�6�8���e�J����_�dTZVfg�&�FW[{?�9f��@lU/��rS�s���ʣ�3V�[$Ri��	oӥE��`���_�I����J�����<�W�PYX��{�L�Y.(v���;U���ll�ޜ���Nw�',�:����P��Ϸ� ��}���4oD)�N����{�җW|̘�.�.���⥵�/�ka�|r���_90����i:������Q:�Q.ͬ�1�XN��3f���h�f��W�a̘t&��E�w6��3���\n�����6�V��r�����:�X|�럂����^��a8s�$:M��'��'J�7AZ�5MI���?��F�h���*�$+�����zG@)x0��0�\�����ޕ�]�v�m��YAy[y�k�D�ӄq������,�j��L7E���ۜ�tX����"���J��?���P�u~�j'��`�����輻�Z�.M��2�h�3-eM�m��g�iT�;�ac�P��/���bpT��
&�&*��V��s%K��p��!�jN���g��?�S��_C_c�M^�L8�VKo��ü=�x�#���wi�����=W��:P��1q���9���
&I�n��#sD�Ӻm��ge�7����ta ��:|T�[1MP e9�d_a�F����� �2�e\�0��;������^-��/�k�%e���/�2�˻���(��5p��ԥUHt?\���ߛ�,����i�{#���r%�s�����+�j��qhN�>��*�7���*1�5>;XZt��@�
�u7X���4����(��?�"my��Xk��M�43�lJ9�h�����r��ؕ��X�E�6D�z�ԑ��w�-���=����W�2*�J��д����@���c ��MI�� *�W-�f���դ���tlȎ��n=8�Q���&��e�śq��z��^"�rg�!��z�?������g�����{}2�yZ�X�r��0t��p�-W54̝*u�3�Hl����u� �x�f�m1�$�^�6���^��Jn��t��k`I�J��,Ҿ!nQ��1��k@�Z�t�<3?_OS%������x��u��l�0� ��K��M�4���Tx1~C��_&�0c�Z�β�8�1@x��K��(�!,�߈h���ot�:�B=2D�;�ʿ�~.�/!}V��3i@ ��D�h�G���US�4�C����7���X�jӼ���z�7	��K�o�?.�q��S%��;<��%�X U�2ü��H-�iB� ɘ���"Q�G�鐓i׎ӏ�n���M� ��Wi��JBk<a�����{t|�Â���왚�b1�&��)RZ�FDF>�ٿ���^��Vʚ٣H���ն��Q.�]�b�.�w�hBLO2�U\Uy��.�ǎ�<=,XQF�ȉ������Q��FX��'����U6���U��AuU�)��6�b%�AXJ�\ �\5�h�ы�*�@������2e���u��7B�o��~T�{,��-m����>�|7��]�0&g��(j��)/���K����i]Mp�Z�O�{~�C����E��pK�.%��	�X���q(���(��
�8?���'V5`*�v~��o����t��j(<��8�q�/��јtaQ��f�!�`�񢄒M�X�˝�Xk�E�?�X��� �5�+����M�٫�|&wf.5��҃��m�/pM)k��{�G�~�ގ����4�y�k�dHT��,�	�J�o��{!*�"
�2|���h��,}]�E��Ƅ��XyJ�j��e�R���f���s�B�B���2���;�"I࿓�]U[�~w��9̚t"r���O���H����qX�Ɯ�s��Xg���^�S��WI��ׄ"y:�(��H��Fl'������;")9^$��� �F�J4��$�H�����6�s'�B��F����=�C^1a��lQ� ~�nŵ��P	�,�
�3���Q�]X�B9�b��j��Լ'��u._Y�Gv�����;�&��xY �mnGÅ]'z]+���������i�"e�$�W�[���s��q�E�����O�!⇱��ؐ��s���c@���1��D��.<�UVIB�gxIo6|����m��
o*��"��I�������/s��	m�^{g�1�nÚ�u������i-Q}�,9BY=���/ާ�NՇ�pA��F�yũX����<i>82�mRޭ��[�������wM��q8Y$��Ӂ=hu�J��7��s���%8���ϐwX�Y� 
�ZJ���ɂ���d��C��}��'}0k<4G,�K$���r�`਽��ۉ2����1(�1�Ȼr�W����]�N���^y3αB@]�Oܟ��>�
g�G������v����M�-�$֡V��؏���Gz��r��x�}:$[�4��@��RU˚�g���
�w(��+5���=I�7��n�ʥDx�  ��ί)��+���OX�_i�Ld�lXU�1���m��� ��(�9\�)����j�0mn-v��7'ݲ��Ǖ� �X�exc*J��g���*���"e����]L�R�B|���F��z�+��w4�Cc������a�����~B���R�S�s�?�@̶=P�n�����Ei{��O�RuHw�~\X�2R̈�i�zO46y����d�>qhy��.ۦ:ޔ�{7L���R�����r1�Ke.��%[@��a�5����sb<M�۾F�F���=D�g�H['Żl$��(�=ͮ�,]%�Q�6~������8���l�<p���X(�M��8u�S�8e �q��<�.QT'
�
�HsZ;�
_-�A&�m=TA��6����'2�.�V9��@�_�@<j�����u�����@M�m�ۛ�#���m(�ªm�t�=ej�Qz�b~!�W�p���̴��/���
��C[�^턃qk��f�/v���@f�M(��@W���pb���;�LɸΣ6ߡ����3Ow��F�,�e�甈(½&$hI������egp�34��e�8����t�����Ӟ]���>���鯫��tG��=�s�`��䣊D��G���3�C�`���T�i�*lh�$�*y=
�Q�YaAvoWY>�@ݻ/z��b_�"@$���P^Z�T���
_���R����.�J��U;�%i�Ҟf$CGq�U�My~V���"���i�h�?ߝ���鼨ߙ~`�#�^P`��扊^�_�8�kQ>�%��)��"-Q����^�h8�ʽ,c�]@��d�ڋ��H��bg��J!�����:��p"�k����Zӷ��pJw�]6���Gr�t�o+w7X״l:,�#�M��R�T��x��}i�}n����p��T�B�\�p�hc���K���_1���H���{@u�l��}t Ϝ��GIM��K��(�̷�z��{ސ�ZiS�:�����������D�"mX(�Bx�(g���pX�h��#>���WR��"x������ES�ƣ33�����n�f��6d]��l|S��Dƍ��+�>f,N�[�\�Ьf�	�R��q/R��u�pޅ�Q�@v�����$|/;���.#�\J��#0\��i��

�b|z~�+���~f�6�@ FͶTc�:M�h"]A�-ɛ�@��[�Vb�2���I|Hf�	v06�\�0��M��A�b(r``���+�8�2�Zw	��(�Ǆ.���/%}C�(����'=�T������;����X���/��/Uޞ5�o;�xP[,җ��4��m�v�|0���D�Y@�Z�<�wyI�~ t4��1,��=�`�ԍ�lvk(�_b~.ШTs$�Y�� ,12���50#vS��Y�.��˔E�����th� f�N�z���h�wSP���@��ܔDH�t�[P��aͫ~S�n��g���覵p|��T�	��'�`3����=����,���/�_6a�zNӀ�jy��J��-�_�[qM�U��*=;��p͵GRN�@�����du{�%e{;63���_1�L���JFd��/��=Iƽ��$1� .;&��G�
�79J��ް�*�#�6y&�D
�{�G�L�̓%�lTlB�'�����Y86�b(jM6���y�8��݁����y�Y:�4��x[5��v�=0Ց8���ʻ�|���5�{�1t���#]%�/�Z{=�B����RUz��H�+Hչ��c��#�c-�1���;�k�#�J��Y�(�A>[��1a�z��[���#^G�P�|m���To��A
4���pֶ��#x0��uj�����\é*��/���o#�!o �^a���
;"$��.1N7s��_+��F)������77u0v�.�v͉_�L'�]�rI�!��(�\�[63՛J�r������"nR7S�1y�w��>luU
��=QVm���T�>�
.��d�Bm#�Epb2F2ŊH��;�?Z	����P6��!w��zI��y ��L<g�����Տ�33�g ����1�pw�����b:�zQ�a���\-��R����:`�}o�	�i�R��\~���no�R��J�}��f���<($]%����$��fs�<ӝM�CQ��[�s�a8b�����[��0HXHtu�;��v��C��7,�]	k��!Oc�h��#:/��O��Vϭ[�m��!a��R�ٰ����k��=9u�߆ )*���-���e�ݴo�ܾ��N�nelmQ�_dC��	�>���E�q��#M����� �`�t�j��0��������Z���bN�$��o$��x͗��F[`� 3���bwp���,�P���^��!���Pr�����̌3V�puA	=�6��lb��i��VQ�� ����OS~n��<)��iu+9+"bMɢ��ĥc�P��k䣘�t4�.8ح ��Z�XK��]�v�����>�(�b���[�W܋�]*,�2@�ąKU�UKH$uA8d��#���d�NO�����0�s*K
�*�/2��	��h�<|���X��]��x ə�
�g�T;Xf�5� ��B�*��
��pXu��n�����w�'��
����0f��^�=>���Zuye?h�=����k���:�<�&�#�ޒVn��z�ֲ�ʞ�\�͋C�$�����8�yt�Z�C������"��*��v�N�,0�0?�@�Y-mT�L�Q�����ʽ�D� �qmU��&� ��DJs�_kٹ���f��.�Ռ�bWGˬ c?/f���C������܃�5�1�2!׮E,R�8:f0sڽ���[O�lB/Tێ&ys=�N��4-a�b�Ǟ��W폈�e�@�?��4Y�=��2ė�:�6����	��JF=���O�9JyW_��Up#C����IA�p�����Uj��I�vf�:Nz��Q7����@��Jp&� `�\w<��G�'���.3x���(��9�U�X�	#�ƍ��&eK�[B��'9�S�8����B��%�\_�@&�8��On�ƓZ�v��+�-߭�&Xry+�Q�k5L���k>m]q�H���"2e~~���'����	P\B��r���p՟v���'��(����>�l������8P��=��P����dZb^��T~0||���ޖ6�����u�)
����_�,4 �r]ժL�7dY� /�JA�X�*���,�}9"ٝm�rd�X~��*�8�7��wv��>������ZYp!D,^f r(���?B���u6U�A2���@�WǠS�ǐhh�<j�1���,�i+(�ګ�5P���a|4�2+�/X1�����q'�6s*�A��:���9#V~"CZ�Z�ϨB!L��.VD�Q���v�!�tx�+e�Q ��KZ���XvǰNT	�����y��:�\O��PS�\�$b�_��`l����zI���ܝ�u%L�M�ZZx,d��Q	�$`ی?/(.b�w���a�r4�MP|r���Vt���|��d�a�;��Wb���5�[�l�J��9�\��uKV�b�F,L�E[�����0�e. �W�`@Y��!�������>����<*`
�!t�}q��_�j��-T���g��:�����y�ա�+�\�}�2��3L�u��]�=q?�f�h�FD�B�]�kv���)�^�]��s�	l쟥;b/�F�j�4��*�y�	G�������,3M�2tüb4����G��#�, ��W"9>� �c'�6�E�M<��/dqŷݽ&9P�����mԞ�t��r�B�4��?e K�Bٴ�ғ��)}9V߰��t�V��R���n$
�A� اgi9@N!�'��],(���J�ci�yG�.ҩ@���b�B�f�DHf�F��A��&<`|]v
%:��:�n]�L���0�(w/cY���Y�����L��H�p]^�>�$.ګ�A���뉉�W����y'`}G�Ym\�|����7���u�#��=�k7�v��;�y��6p�0�޺���X�*]��ʛ��Gn��A���2�4BS��6Y��E�.���;�0+�/x
i��F2Z�����t���|r�[ԴǕ�i���/�1�߮x�����#�n���7r������ӗ3�|޷�-��t�q	(\���f-#MGj��|O���pxw��7�ѯ��ASl��vn����oBLV���N�m�Z�ה����	��ķt\���`kX��d����as��,~_��cJ[C�v��xKoɸ΋��cEqY"&Ρ�CD��q�3�8Y2So89 ���V�'�R`9�/�Q��9E�=�uʰ��P��:�9�ñ-�G*?�~%�y��HJH��k���Σ��qȮ?�pZQ�~ɻ��,��l���.��S��5������2b�w�~9e�}'�:�*5Y����f��I+w@�[d�� �@y���҂R����i��v
��=��>�#�~�S���%���+��X\iI�K�a��e,H�j�X�O~�0�=��c�U���B�*?�I-����zy�k��R�@�I����)�2�7oL�A�z��k'spGp��=^��m�{J����l ,(��V�/��s�"�z��ܛ+�WG4���a���uߐ��b��ako�l>IOMiI9"�5��B(�?�V�|T3n�]{S��>�ֳ��r]�A��ҟ���%j�����E�D%|Cn�٭S��!����'C-Җ��u��U�B̠��)#�x�F��v��⃆�Y�*�鹰c'�������{�o�h�8�pD<E�A�a�������q�r�9�'Y�g��ھU<׶N�wd�iǨ0�|0��ϩ@�[3i��!pE�� �Y�Gl�$[�1A�J����'���ܺ	�GY\��YS��+t���{h�~�Y�aEfBps�VhM^BZ�L�[�@�_�5�P��BT���G����rx�W��c�~쑾�QL%g����"��wq�?iL3'[&�E��b�	kgle�FB�9�3�����u����+���N�bd�i:%��p����h,b�,p���u�_��مj}���;4`�X�� SxI�](#tN#��^��=�ʊq�Z��;���(�T
? j-��6
�����-@r�Q�^�Ō&!�͉�5��XS@c���?{DSW�ӕY�}2֬ρy2�����w��E4��\��	�<
Ȭbje��O)y��5@�>���z9��ݥ�xx����n�*�윞�nJ<ռf�1iVPϐ�0Z_�S5~�0��8����n�o�H�_��5���,N�L�L���y���rr�k_�T7���wLH��,��|�3��n��MH��9
bCV�y��� �'L��L��;�<�NȎ��I���җL/a7ZO����ʽ@#MYJ�C*�֖M<�owp�	bn�v����
 �ڦC�e% 03�)��Я�K<����= `��H���\��dm)����؏FLb�f��Z^2��O�zJ�'X�L"��h��K�-��H��_���i�g<V��O� f�杄Uv914([�Ԛ��ǰ�F��R!�2A�$�!�ګp�ƼOf�73������Ug�`��a$2�c�'���F��7⨵�*L��[x�ё�_�����\4aҧص���KZܕ	j�|/h�
�1�J8�5_�'�Z'�n�z�^�/��*A=Dv۟�-�t'���c�+���o�0]�L��do�e�(��{�E˵��uU%���xG���+[��Vg���^�h(�
k�o�=cT��_l!0��c��7�C�L��'��&�",H�-:���c8�Q�������$|10)\�G�I JY��#�aE��+��[8]���.��o���Y��
L(�x�S��}�c�ￂg[�H�A� ���+��@���rg&+�U7"�?z��w��>�c���9+A܄��a@U z��ŠᕢE�����A�p�o�1�H��X�`xb(��S�˾:������8��[�L=�evϦ�,{vI/2Z�zO҇���<btF0�w�bv��h
�7'���;�l�{r�L;� [mlҹ�������}I�k�Iik��'x�~����6��ʝ�T����_�5���N�Q4$<<�J�<0L�N�4m3)��jE���E���C��y��k��FDr�Y6�W1Ș���5��i�K�C5�����������
/��M�������҆�ɗ�R��b����
������d$y<14��RK���>c{���Ix����3�7�&����ܘ:����&�����٨����a�:jc�I�w��:f�?|F̨�U�/7�xc~���D�#nB����6��%_G�Ql���os�:��$5�Aъ4�D��غ"Pެ��}��&��L�_�O<�q�O�_��͞|^븎&iL���Tٗp~7���9;;�y�G����i�����*���x��$:�@|3ə�. K�P��s�7�ܛ��+6[5��_H�Z7�*��j.��Q@�D]%�]jA��S�
���)G��E&�9o�3f���vP%�e3sv�w�����Dyېi	zȣb\�,?P[��d��ƚ��<��4&QB�8����@��5�9^�WdL{���Ҩo��eP���t]Z'=˯�̶(�P��8-ӞG��$�������S�8�{����	�I�w�jD�g`D�O?����A���M.3��)]4M������J�J��V	��q��"&&�w��d�=PXP}�;�,��p��������ZǇqZ�7��(?2�]���t���v9@
�֭�/�s�x#����C���Cuj~z��e�>�Su��l�o���)����f�~Wj<N�X~�6���W��������F5�%2E�!Ó��&<]�<'_�\B�JM !rZě�qv�0K��[fm3���&�����
��â�HD(B��5RK�2���Q#���P�s4t�ZkFr]s3l�-8�5�%��EQ�p����J�����4��(SCg��:�Q]��h_YR���<}���跲P�yAC<B��߾Ă�?:��)�Ș��R3�,� \�u8G"�#v��MGDӖ=)��R���?#W�f�/hH���lO#��(fB����
�F�8��n���ф�D�	���w���ˁ=���Dj��UUlݧ�y}}�e�Q>�%"������~֮��(����G�Xl��Z��
�l7�Tê۲I\'�#W�/���Z
��#�9�{���
�k�7e���Q:�3�q�����w���%bS3�y���>�����9_���4׹&���t�֜�T�#
����(��ϟ��d�3Hu�2L�aJ�u^�x �����Gл��Z�G��-p[RX��uv��Z�� 6塭�. �R�[��b�I��	���&/���ޥs�������Ƒ`�6DMC��ر�t�� c����[���k�H�Ӷ����ޫ/R��B�L1�n��Dh1%pD��)ԯPe%��E^:Q~�Yi���d��qK��;G�8n&�*{��3�Ug}�e�u_�%&�	Xz=�jb;���)a�9G8���b@�v~"�" o�.�\�&Q�0�D�e��>�����m�0e��Q<�g+��R0/�/�%i��DÌ�e�����?��q &e�Ȳ��a<N��\P��`�'�?��.�V��Ô��h�AR�Ċ��'�0�a2U��d��b~�ꋷxؔ[E�.��I��F'DW!{��Jq�$�f�b���q~=q'^�Bc��*�j��?FڍzZ��$U!-����:��_�̂���K��a�ti@�MR���Y\}&�0�"6'Qᜆ��8�JG߲Sk �t�q���ǟT����P�ı�.D0&�Ɛ���Z�F���P�|��v6� X��1�2��/b�,���?cA� �{W�0>�R ���@����}�H �ŕ�Q��d�7qQx�tًEY�=W�vr*�,��e�ETz��G�r��AK�G�R
[��2꬀eE�<���-�E�W�A��{� 8B�7��ȰUP�gz������q��R�t|���]�{/���V'=,�p��ƒ����[�.2F#�M�b��RDa�Q��E��ō�\J�Q9�--''�,׸�{s
�� ��Ѝ�@��V���ș�Hb9�P�v˷���w�gp�aڶ�Y��r��\���E��O�r�A'�O?��EW����h(���v���Ȏ*�9]���L4��0�Tk)w����@�ӊ�2�o>�/ 	%�!�Y�y��'	S��m�����T��ɺ=+˺���C�[Cq�a�G^D~9b���7b%xƒ�p?Ecr�zy��������_����D>C*��oC��+`Zʩ�B릆\�
����0v�j�}�5��N��	�X^,�DZpn��6)���:W㑓�V�i�z�;���C���)QM��?X��N3 �ӫ�x4ZHo�?��3[�N��w�s俬��7)0*��Ԧ���� �x)�m��( �v��t���ی~��Rи6W�O:ֵoѧO�2��,sd���#���^���rAYS0��* �� 
#��傋�����d�VR��MFN�xkMh%��7|�%yI�k�Xl��:�[�Sq�ӧn�h�f�ٶ$ާ��4��(�c�`�[u�xW�J�p�|�.0Fް��@j�
|3*9F��\����;=aǏ+��9���
ew�Ăg:V�!��jҭ=�C�2�i��C�뿛��N��Ǖ�0c�
,���ސ�B-�w�ߣ��j(�%7eeh�(��xA.���,��k�Rc3_�d"}�m.Y�t-���َ ��1��_­��sR�B�K9����Ue,5����E}��%o�.Q�f�째�>(>H���J����L����#���~3�t� �g ���P8�U�F�d���� ջ��7ͭU�K5I��H����@�T�����io7��$�Ж�:��^c�3�NZ�U�h ��/�`���|8�܆���K��	���pAV�_�M{g/tJFO+3�w�%���]1�0K�Dd�r`θ|�U�FZ�[q�c�"�YH�JK��	䊮�#�=ÕP�I�������udo<�������	(HQ5B�ф�%Z�ٴsA�԰��F���~����:�����a4;�h�ڷ�í���c����+WE/��B���Q٥=E'�#��6d��u+�X\�+5��0�����^�}W��~#��c�+=�to��4љ���jŐC2���*B3z�9��U+�wd�#Vp	����C�Y��*�i (/�5e��hZF�d�{���ގ��E]T�UFY�Lq��I��ѕ�Fd�F4g��+���:qPD�ZZjI#�ǜs��Ùu�7�Zq�@��$L	�W&�ʠ8�F�~V�N9�w[���8$;�T��*�;�<t:�a�@���,���*��C	�����Ɲ��"�'�z��_in��h�6w/�aXyￄAs��<!�ʑ3{=�#�1�4"m/�Ϻ�|�Ĥn����m�1�k6Ga�����5`$0zT�<��_~NH�+��{���un����Ÿݯ��H*usddl����[z�]�0(ђi����x�w~h���K5�KobÆ{��1��}�Q��!I�o���{.~#&�6��'1|�'�۞�s�Nf��3��D<17ɀ)Z�}�=+k?�,ll{�Ӭ�i��/:& �H�j�S\��Ʌ�Iy��ŌDx���5�!ݭO�{��Yk̓Li"N1[Y�seX���S
�({.���v�ܥ-9uɤ�<$�<��'&���dr��˅c�Y��˳�/Y��T��`��N,�~:z�N*�͔�a�l���q\��Iz�)��}T²t�t->�~H��	j�g�cTL�d�JMHz�g�	�NS<Ή�V�����hſz����<�k�%g�E���/5z�ح=Cs�1�l�/I���ya�#�����2���Z�Bt ��W�i�K:�uř�c�E�Z�4ǖ�)e��r6k��5C&qOrw��7v�����WS*��]�P)������@7OMR�/�	��ZN��/ Ce>�a�f3��+lZ��y���K�.�/�g��r��x�^T�l�7���v2%=`-�OV���h��9_g�]9�a� :�WSL���K@�)�<CsW1�����N�o�O�~�}*�	j3=��(5Rń��r��;h¡��LB�C�+��ҿO�Q2�����N��)܄��h����{e���њ�g��aS�Q�$�GG|{νٞ4 s��R�x�F��DP��4q0���Gjl�=������r��8��BIqu�؋V1w�s�&�i��6�}VZ�!�S&=��E;���nD���4�C�ڤ���){�����=܆�iB����v�{�F@�ٻ���0d<<�n��<pH��	����O��0%���۱�x���١���?�O����^�r�9ζ����^G����K!�r��KƸ�%��!�Q%D�_�c�S��ke��##�ӥ���`�2�0����EZ<v=ۆ�<}%&g���	��p;T�&!7H���uF�@Tyغ���l!Sܳ�`���g�qZܮP�N�7D������f*��"}�*U}+��d�P?��<=�Q�)g����7�x$!<�������`�Y���@ΉI��C�w�7i���?���ƚVM*MdzX���s���=?y�Yc�/��eR�;�b�{A��Q��T�G��a����V��.|T�r�$˯˳�Ȱ��]ۼ��\C�g֓$�zt����n����R���c�'�������0�M���Wi�����#Ѳ�|�6�n���B�N@�<��µ��*;�k�@ui�M�������QCL68gr��9���<���9o�`�x�	�E�W
V<K'"79Լ���d;��ڝ�r�T҉̔AЏwk�4��^|�����}���8�!����f�3f���R�l�/��'U2��?0����$��F���6]����-0�,�":sk����r�:M�����J��f�Ȣ�y��B��|��4��ͽ��ٌ�)T��S���x�}r���������x��)0ҔC��պo�����-͑+?�
X9�����hioꋟM�?Ϙ�N�9DO��E����R�n��������I�Қ!	�>��^��Oэ�y��˵�ؖг�e�ÊCh�_���>���nr�}X�y�_�1ʾ�\���3����е�^z+4_�N���J-j���	�	mϗl՝}5V�!$�I���I�uT�����E�u˛H+����?�`��W45O�:��N�ts�0�}ߊx��q����<@��)��Q;����д*~F��lc
��<� DNlvJP/\�K�����ǫܯ�-3L�ڋI�	�>@IL���NG�y3<2�}� f�5�`�KAG�#H����X�;�I����Y�m�f��RvrH��T��;��i�y��.gY�&c� yT�U��I]P�E�7��8��	.�Y�-����?~���� p�mX�H�86�|6h��_�sz[��r�R�w����2r�'�;y"�
���.^!dR���1�'��89�^�����1,�OC�^�p�I'��w�p�qS�$TQ�@���`�v�Ef:��E�q�����3}�]��SnK��u�`�Y&<�� ��3�W-��ܙ��#�$�e���F_*�f����f���&�_^8\�SP� �W�p��6����.���uw�Y�`_����_����8�`��{��ן�n�aL#z�zD$Zfh�YW5�+G]4SE�FSa�V.2K�h�;�b�
��HJ�t�r��>ɵt?� �_p9���'v�U<��b��������Աl��c�N��&U�5�LCD�#nB��ܐ ��	GT�>���U��^G
��O)�'@P�$�-J=�l��ט� ��3ZT�gEg}F�Ϙ!��� v�s���c��ΉP���O:ܼA�o�P$�mOSMK���7���x��"G;��qZ���¨����=�����$��rb���@!DE�nl�\�B��(��B��p��	QJx^c+�Ǘ��<�v�Lihc��_�]/�5~�nC(]�t��u.�v�5ðx�4���c@�fnە���S+0G�B�95g�bU����*�~��8��*1�i���qw�k�B����0V�ס~��#x��\4�e�(`*��D�+u���6��
>�R�� A�j�_�x�!
SCl��1���nG��\���U�A�����9�.S�QL�62�Ҕ� ��,��***'�CޓT���&>;���/��Õ�/6��[[�ǗB���O2�g�:TQH�{8|�~e[�:&���h\H��q����Œ:�'x��D���:���n��i@��1�V�Yz��TG �cX�H�i|��gV٣ع���G���Q��>�Q�cq�wR��'�չ:0o~�S��p�x�������0ȡRս�5�eE��q�yf�`�QZy6a�J`��
�!s"^=^�j��t��B�e��i�8F�4�{�YZ�_�U'ǥ��T�U2���p�?�S�2\�{KSh�����j ��.��bl�,���B7���~���b�u#�6�)��	�JV���Eڱ<��!��x��s�n��5�L�k�X����Tg��|$��n���e�����L�J/�HY��&֘.�)0�9l�D�I�Y��Q�^�Y�n�Ș�e/�^�-J����f`>}��ýC�Bz���A�t/�@�{X��L����p���ye8x~Jd<���8��`�n�)�$b5�Y�Vd�yw깰*����$N�w�{D:�n�g�xe�M�h�}Ufw��<I�9�(<ܨ�:���Ee��E)��܊M����-�&���[^N�ȿ���E�0yME��ץy���c�'h������~�r�����yO`H��E�������o����o����kE��L��}.�kKb������ʴ�ұ.��w?
hE��
%#{t}�[q�;�?e�:7�9gmSY���P��RQ��g�^�LN-V��A��}U\�i���z�B�i�!��涂(��.�0'T#��wZђ�f# HXx]m����ŵ[�T��S�#\�������P~`�/ݺi0C�|9rL[m���)I�b���5�갰4���2��։�̜)&��Ld&���j),�/s�>[��"���wpA�5��H�y(��k�	�V睴7���H�)p9���Bok�o!�e��6��a���Y��L� J�&���="~[����JG�1�E���=N��ʳf����
���X�^�q�����.T)w�N=��|���K�$A�E`<JS���J��q��P@ w���]x� �#F��^�D��5}%��e2a�4�����Ÿ�υ^V/a8�����Z����k�4G O3~�����ν��y!-ب�����Ni����j�H���atܿ�:�f<+Ƅ�K[�<P����<	� ԣ��R�����U�/�����4��}e��|»�0c�ͦ�¦܁���KFtMT��[S��S���`���)(��:e��%�gH2G��<40�2���Wj�¨��|�`�-���nD4%hZ:~3���(�����7xf��c�(�+�K �ȣT���A3�������ǫӖ1"N�c@�/�j�߇��`�[ݛ��=�;Y�xVZ�E�T�h
�?�~��0x^B$�̏�� .h�{��֓�݆GD��֊��+>��/��sSy�=[�1�+
z��N�	�^��t�`��s��Qg�����޵+A��C0�+�5�)v�s*�1���{[�4���^�\;a���΂Ƃ��5�B@�)�7޺��@M���I����FG�א��G�FͤR�
7��%�]�RC�%��މG�S�Mr|��- 3ں�U��\�(.����>~}(�B5e4a�t�.�W�?�&H_�c�c��-��P?�!٤�eo� 0���Ē9f(��)��3i���)�J(c#�w����R�7��ōھC�mR�$��|�i��)��>�*�Z;=,%�4زO/��R@]$�s�X�ˬT�e)R�����ؠռZ�j0�0#�$���i�2����.>�d'!:���)P�N���(��e|� ������X�	H��d�T�˩y�t��E-��;��`kn2_��k.Ѝ�h��ڽ�O�E�0�	m��G��u��PP�4,��	y%�bK�k���;
G?~*��3W��D�M�|�qy�,&�x�:�Xܹ>/+��oO T
;�Zgr���4=S:��L��p�g%�2,����y�U8�~sjVJ�k\o6�n�o�R^��>�X#��iwO��N�-���cB����~3�� y�Z	���h�� ���4fo7����U��V1L;�	_�d�Z�₝޳��t��U�o{��* P�q��n�DŅ\�͌VHN�K�Qx����GZg@�=�u��&�XK�n��T�H?�ĪQ�^���Ek��6��E�aH^�������јlCW����I�װ��~�X�y����T�o�����NI{XE�n�V���X?4�A������0L〨!�P.us�m=��<�GH��-�B���`p1f�64h�L��h�ܩ�t�	��h����8tݓ�!�(j�<�h�u�r�!S>�ŵ��y] �ͫ��
;\"���s돽��"э�pv�\'��d���Τ>OP��O�X:�= �$`O�8	8!~v6�o;9�-˹ٚi�i����C�ju��{�?ChF;���Ǥʇ}8���h� 9q���(��{D�j�����UU3����x�l�v:?��;%Et��>�(��$<�����M7�9:�=<׬ߓ� R�F�m�x\��Ƌ�QĤ�r�b�t46=�r҇BR0m�5;�f#��"
u�*���i��0@o,�Xt�y$�񮑵p@�D���3m�_꼣#�!I0��)=T!`⛾�
y���D+���"�\K���s����Ч��)G �
�Y��і��������Z�^��緈�.f���\,����׃�\���&58vg��L��Xr��{��aa�l�3��0R�b��XO��f�ޝT��@���~����`��uǰ��4.�^b����Y���A�*�D{��n�$f
%��E�ģ��SY6��	�T�+���>�aٖ�,t���t����1��|d-��⎎0jGյ�g+,ְ�.� zlG`�S�ت����H��-�U���hec������mV���A<��j��65\��{1~̓��b�ĕ�szP�C �V?
�~�& �a����{)p8��x$ ��*vhy�n���693��1h�s��(�;c�g��F̵���w�����Z�jZNrP����s����J�(�p���?�Z���N�ʓ>내U#��;��˧�M:K]00���F��!�枙�\'�n���蓩�N1�S����eRm�^]�$��7��$ �������ʇ�ږ�cLn!0=��'P�
����,�嗡�v�zC��m��0�7�x�uŠM=�1���>�3��0�Yч	� .Ŵ0'�"\HA����td�
�^�}Տ,<)���2��~���������2��N7�_�:B<���ܪs髜�~!k�#��㩫R�"Z �]�;��"��Xx�	(PzՋ�]@'M�r1�U�O��_��dͱ(�Y��Й�~bøOEM�o�F=&�(���$=�:�yI�F�iu:��FZ`�,�;l��?�{N���~x���I
���R�]4���MDc�$˂���o�s�ŵ
(��ͽ��ph�L�A�kґ������tF����n��}e3���� G��}��Q�~Tw؝��\��$�t�����3FTf�j:n/Ij+���������T6�-?��/�m(�V�7n�Gz�K���Y}9Ol6}�\	~�J`��?T;M��|��@{H���6��۰"��꧶\?��)��J��_�N����CH�$�2�iT"�	��2�b�"��4`QT�j茢p�?Nl �%սx��-���v̘�=���3)IV	J��1�%Z�n;�C��&II��9��Z7T�����-@�C�vU8q��t&��8qj%���IL��س�YB�Rt{�\olG ��-���lz�����+n���T���͓?��2��8x#�������֊��DF#zt޸��*a�rE�I�e��~,5%S�߱wS�qY��_\�����:wJ�:�h�#��b����BDM6N}Q��m7��0���N���>��C���Z�Yt+� �
b�!5��|�0��^�iV̉j��ݟ�Q�㼤2ڞ�@R:(g=���/��'�~�D�f-{��^=/�>��(pFg>�1����@�T��|6E��}��d1�(֔���G�����6u&�P�K�qm��ܖ��Lu�y+np�.S�'�\�<�!��^�w'�Hu���^��4�Űo�[��j�AѰ���]���4�V�Lcʊ����jwl�@�PI�ݗٺC���}x�y��[>�Ƌ���Ui~�A�6⍚1��cץqo�:sL�����Q)�������r(+��(�:������/=S�Yf�徕�O;�E��VW8�W\�:��tM��bFv����cY�k���f����,r>��N��^���xa�e��$�Ȯ�y�T���R������vF�#^l9d��1�
㱡UE�,�I�k6E9����+�;�nON(VdT~th��d�R���Ix
�'���O.�J�q�~�=����A[r��Ϭ?��n���S=��2�f��~n�ĶN٬�G&�E7��i�������M�)�vn���N���7M��J����a�un@4���[�i4NNk�{������3?�WH�I����UL<ڿ��j�eQ���se���@��ȯl'1,��)�r�M�8FW@F]j����5�]������cl������Du�s�^ɮ�yP�s��T��+���e�ES-��������X9Pʔ}�H�@o�
�Q Lݢ+�&��49��KH�=�|?��r(�`[%8��1Ɣ���F˳c�aW�q���1B�U�l����Ȗ���4�ܙ�'Ƌ�t�@�Шfhf��<\`�}"�ѐ��!;��4�9���TM���Y� 8��0[��B�搧�s~yI�.hx����n�N$�ǶK��h3��`x�;�4����;��a�^ʕ�)9�Â��6�����U���F�+���5O�"�4? p	J�8NOhL� ���e�ļ?��k�3߲rL�^s��w��_����+���i�W�䣩?��yF�V6}�lu_��'>|R�<k#��5���)�d+�(��������ٞk�b�֬o������q�Q(M,⸊�oЀ�6��n�~z���Q�md���B���P�C�i���㢛�ky&wj҆��(��㭍�̕i��P����a�&_��Xw��+��6>KaP�C�c�5����*��G�&X���A*�;��U怳)ly �Ǻ�U�0���#��ܛA�8:k���^P�Q��"F-=��z��;���8W~2�5��L%�M� �Ot�~
Q���䖏�o���mN�m���	\��ty�'o�؃�QJ`��R���&��|g�c�x�9��LI�N���V%��w��t������.���Z7�\�}Z����dp����A`^[���K�D�y�̙�Y��v�/O�g.���4��כ>	��PgZ����^bcY	i���~��ͺɾ�KM���{��������Ɛ�΍�8y�:�!�7�V���ݖ��Τ6k5���Z�X�M��Pw�V+�t2�A8��l���X5΀�"3%.[�0�z->�J��c](<�E*˵V��i���:'���	F'�vĵd,
R�ө�4����Z�T���R0����Ȱ���r������[� R��O����6<�����[�o8J��1YԤ��Ets��R�2k1�J����}�|a\�`���4%�K�$�YJ��q�u���Ɵ���CDCkC�9�vֹV����ԛ�W��؄��#�j�*�I���D�lWف��f7?p-��H=+n�{�qqO|�p��4��#1F%"p�B��Z����AA��,���nE�Ѡ�6Λ���Gz����.nȆc;J��x��R5ڱIJ�=mU�~�Qޏ<���v2o��gs�l������C`�ݴYS���Ol��6\��'����Ua�b/!�W+���x���5j�p5N���k���9�Fqʑ���?Q6E��nݶ���϶�4���+�j�:���>�Q�o��r��Lz�:e��^����UW4��A�f��`χ�6@�%����J 1������ JGR��,��ܚ	4�����C��e�)T��/kd�ƕ���f��w���Rx�;��).u��p8�֣1a��)�%^��Z
�橢̥�s��;�?dH�����5諰�������o�N�(���3!���F���܂p�i�G���|�����)�2F����Wq0�`۹�Q�*滉]8ȿ���3��K��'g }v ��;+�T�vI]BT�%�YQ�����R�������@OD����5/Q�Z�	qx�
��c}]k�̴+�:3MIg�2)�s�xk�) ͥ�NW�g���u
��O!�_���wW4��eH�M�[1�%�ֈ����˙k�������fwZ��A��Y��ꏺ
�.���qw���
u�x1��k}ۧq�>�hk�����k�b�Q`}SB��'@r�u�v��C)
�#�I��a�Nl���=Ȕ��ƨm����;T̉���H� �8Ӻ^���5��Im7��JX�ƌ��ke��a!���fg O��!9�f��r������B���"y�G��W��<�%���nZ*^�ej�At�[����gb>=��*�!�/VĚwC��lQ�4�b�#��3��.
��`���Q3����� h5��劽3��$�<w={>��L+p�M�x(��3�E�j?٩a�g�zsҮ�8#��J�O�+� ߄D��p*s��3�[�<�mE^�� P.6C�ʨ\�&�l�\Z	`r��+f$��]���m^Qʨ�z���B���l�̋ՊO����xo ��4�1���|b�B�NM��F�g���80�9�.�&�9x����-�&���1.J�������>`��e�L��ٷ��?���w�Ja�
�\Y~"��)��R�ΘK��R�Mr@�(0�-ӳk���Z�]�󞋍�X���U�E�]�>{<)4C�˫�������rB��砕��q;L�*	�~hp(|�	�l�RC�Y���>oT�>��)���.�R/�{�s�5pz�B��]����;v�؄3�p��M�z�
F��B��O���%(�3��`���_������M�K��
�V�D^5p�Ý���H�	AX摨 ȶ�pR�1����@>ƭ)��GF���?R���G��_��zm6�~#i�9l[7mܙ0cF����bѼ�g���{P4���[һ�t	Z#��F�F҂��K�g'q|����s �x�VԵ劫�ӧ�o�k����E���p�ԓ��Ҫ��w}�,�+��) �h�M��Q%��H[+}��f:�IU�
�-�|��E�֛CM^���\u���L��138�ܳQ}�f.'(�`1�xmЩt�nhQ��w�_Zp�dӫ��3���-ǵ�w�s��bVw�:l�p�:��?��䔥b�w��(�����a��{آ��l��+U�u���6��.��G�WumO������d��I�w�6�\�_[[m�Ҥ� i��@P�Q�JI�!]�^���}6efv=��^�y�~�Gc��8����Y�W�Y�i|j�fg�E0�7�=�(c�]�\U���F8p����o��V������ޘ�\K�"9[&��R���6=�ۙGx݀�e �fyL���d-�NK��t��Г\??�:��5ZӦu�����;�P6��) k��W�#��N[0Λq[�C�S�Z����������	�b+�)�a8�Y�ړ��]�09��R�iT|��ꄅ�J|
g���m����r�uU/Yv�C[��W���O&�=Յ��4�Q��z�HA��IO�iE{(���ҋ�+�i}��2:�ӉS��t���o��?[�t�P�J^?E�Df �a-�؂W������\Mbd�4�ל��j|�|�*6Ȝ.�w?��Z�Ff�3�I��"2num�A�@��(Dư�q�e
7bΙ�22��.�[j�y�J\�Yb�� +�~�4�hoȴ��X)��]Ȋ I���QQ��i��G���N�ס�w>��SS5P{��||s5T}Ǒ�K��tn�`���I���w��+�C���W��1�+�r�YAL�ß�\L����("Rji_�JЉ�Qf}?
Aw���H�Iаҥ&�HH�hI/�tp,3%��x��"��	�;�#�T@$���n�_���8�ٺY�w\�%Fy�9[�g' �J-Z�e��Ư.9��"�4��%�ݞ-$I���ul�KaC��0�ͧ*钂O,V�/Zb�/��v@�,@%�c�k�S���H�w�F�5�8#j(#$@7n�n����¸�w�bT�g)�.���`%oA�l�a��e�����gʹ�өE��j��B_�B/--��z�`�j!���|#��,ppC9n��A�k�7*�A��u4c?[ড়��c�>���v�
Mȧ���؀nT���s~(ͦD��P݉�}�UAm��w0�bߍy��\��m۱,2��m��Jm�+y$I�[�Y��q���>���[E7�{_x0`i3�j0$%(G�{r�X��9�_v�t.�9���5�N�R���bA����<����� /�E���R9���~���Y�Q���v�aKq�S\+S�-��+{#5�:���`�4A�N��2���q��~V4b�FS��*�, ��ɋ8�˻��/��e�����rC�NO�W�6u��C�pQ�ɹ}M��G������H8<$lو��=��$�T+�}q�D5�����*��@l��o5oSȃ�4<f���� �K��%d��� �%o�C��lo��"o�^�`�h����<.��z♇�߭��|��@�FRe��',�t[]���<|�OH���^~$7�E��
�U;{��&X:nF�y�ǥ�)����¡g7s���\ѿZ�L�V�A�u�M)Z\%z��I�s�����ث���t�Wۖ>kR��:��9�n��h��;uTqR�C����Lc(G֢����RFG��C�A_�\�L�y��9��b�>V���y	�h��*7�?��>yi�'�ܾF�S��Yr�M�Z����4�݆��h�q�{��/��C!��.�&� ����zg��dާ:�qh�sO�%�~�+��'�ũٰqB����#0�z7�j��!ٸ�#Ж`m�R� Y��Jbւc�+P2�m B��W���[�)]�+�$>���J�&kJ+����a��h��58�#H��'[� �'��Y_^l���K��L�`�����|�CZ'��SՊL\i�\��Rxs�����D��N�}/��e�JYk�W�����~��*#����g�x�� �M��e�I_#����8	A#?�5�]�L~�t���f7�Ua/�H�}e������x���"Ѹy�5{���0)��T��������ڷ�s��`��I8փ�Rx�ոf�O]+��d�u�mu�0�L��T���y���Ӳ
�ZY$՚����Vpy��,%�-egY^���t�bw`���@	�o�W��\�nin�	m���:�@ں��{sWe4=#�L+#��a�;.O��ވ�ꙁ��yŎ�a8H�(�1�5���|��R�m�e7�
J��O���.�mj��i�jAc�3������1��1��A����GU��n�����^=+��{j'��ÿ�|�$���-�R�Y3
�.W�O�.�W�v� ]����@1})�g`	2
c_��2HgC]v�Ԗ�@����b�b����.9.����P˛ݸw��O��c�բ�="z�c���HS�m��UX߷����ث�<cC��auN�y.I�j�%&h�3�������{pZ��ay� �]���r�D����3YڅN;�SwS�o�>L�='`!�3kRԓ)�CI��т����ac�Y���A\�F>�dpZ?(4&A	�.:[_pV�@��c�\n�������]�����q�K(kB��EC���w_h7-m1�5�XR�S��t�>�o�@����g���]�e�+蟮��SM�(����1q�=��f6dK#�S��<M��p1�ԍ�с:��C�8N&�o��2E�E�P�f �s���U4������H����9�.��1E�O�\0O̝���?��L�������$�(-�&蛊��ݓ�zV��^����%nnI�cu�^��t� �f���cr�Y�\�R�+e��4��^-Jq��k����������;�@�����}bǅO��qE".�{�f&|�ܯ)��͵Z��n9��P��:}�������Q��f
���
e�c�b��Hk�������w�~���<�tv������_\`�Ϡ�9�zo���*"\�i��I!\����5'�}�%ǯ�Q ��������Ϧ�%���������I����k_�����f�x
;⻔�\�<>(yx�iz�M7����� Z���:�R��e��м%6g�C��������x��R����u'o��?����1��m�P���ʉ����iH9��r%<������ڜ�<��	\u� )����kͥ푣ZI�]�G/Ψ����r����dI�[P���cF�����0:l�[�gձ$E��&�j�)�c#���KU��<6)�-��N��I�uM�Ӟ�H�k\�3v��P�m�ed�o�"��\џ�	�������tb{�Ba�R��21B��iP�}�07)��1��4�N~��C-`~Z�^���jO~Y�C�x��g��2�w���K1���?�j�J��;4��LL�E�
=�?(ܛ[��b{�\?��uDC�W7�;��`������RW8}�dF�Q�ڜ�-ۤHa�1������~��V���֦�#�����olC{C� �D��5�M0�KU~�����#Ç@��vM